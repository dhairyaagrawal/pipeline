// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 64-Bit"
// VERSION "Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"

// DATE "09/16/2018 22:56:05"

// 
// Device: Altera EP4CE115F29C8 Package FBGA780
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module system (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	CLK,
	nRST,
	\syif.halt ,
	\syif.load ,
	\syif.addr ,
	\syif.store ,
	\syif.REN ,
	\syif.WEN ,
	\syif.tbCTRL );
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	CLK;
input 	nRST;
output 	\syif.halt ;
output 	[31:0] \syif.load ;
input 	[31:0] \syif.addr ;
input 	[31:0] \syif.store ;
input 	\syif.REN ;
input 	\syif.WEN ;
input 	\syif.tbCTRL ;

// Design Ports Information
// syif.halt	=>  Location: PIN_AD15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[0]	=>  Location: PIN_AH17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[1]	=>  Location: PIN_F18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[2]	=>  Location: PIN_D13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[3]	=>  Location: PIN_G13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[4]	=>  Location: PIN_AF16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[5]	=>  Location: PIN_H15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[6]	=>  Location: PIN_H21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[7]	=>  Location: PIN_P1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[8]	=>  Location: PIN_AE15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[9]	=>  Location: PIN_C14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[10]	=>  Location: PIN_AB15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[11]	=>  Location: PIN_AA16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[12]	=>  Location: PIN_AE16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[13]	=>  Location: PIN_E17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[14]	=>  Location: PIN_H13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[15]	=>  Location: PIN_J19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[16]	=>  Location: PIN_AA14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[17]	=>  Location: PIN_R25,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[18]	=>  Location: PIN_AA13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[19]	=>  Location: PIN_C13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[20]	=>  Location: PIN_Y15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[21]	=>  Location: PIN_M23,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[22]	=>  Location: PIN_R7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[23]	=>  Location: PIN_AH12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[24]	=>  Location: PIN_R3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[25]	=>  Location: PIN_AD12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[26]	=>  Location: PIN_AC14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[27]	=>  Location: PIN_AG12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[28]	=>  Location: PIN_J12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[29]	=>  Location: PIN_AD11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[30]	=>  Location: PIN_Y14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[31]	=>  Location: PIN_AB14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.tbCTRL	=>  Location: PIN_AG15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[1]	=>  Location: PIN_AH15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[0]	=>  Location: PIN_AH19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[3]	=>  Location: PIN_E15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[2]	=>  Location: PIN_T26,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[5]	=>  Location: PIN_G15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[4]	=>  Location: PIN_C16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[7]	=>  Location: PIN_A17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[6]	=>  Location: PIN_H16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[9]	=>  Location: PIN_AA15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[8]	=>  Location: PIN_AE17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[11]	=>  Location: PIN_T3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[10]	=>  Location: PIN_C15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[13]	=>  Location: PIN_R23,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[12]	=>  Location: PIN_Y12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[15]	=>  Location: PIN_D14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[14]	=>  Location: PIN_AC15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[17]	=>  Location: PIN_G18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[16]	=>  Location: PIN_J17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[19]	=>  Location: PIN_R21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[18]	=>  Location: PIN_D15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[21]	=>  Location: PIN_AF15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[20]	=>  Location: PIN_R22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[23]	=>  Location: PIN_B17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[22]	=>  Location: PIN_H17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[25]	=>  Location: PIN_C12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[24]	=>  Location: PIN_AC11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[27]	=>  Location: PIN_A18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[26]	=>  Location: PIN_F17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[29]	=>  Location: PIN_J15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[28]	=>  Location: PIN_G16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[31]	=>  Location: PIN_D12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[30]	=>  Location: PIN_R26,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.WEN	=>  Location: PIN_R27,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.REN	=>  Location: PIN_P21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// nRST	=>  Location: PIN_Y2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// CLK	=>  Location: PIN_J1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[0]	=>  Location: PIN_D16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[1]	=>  Location: PIN_AB16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[2]	=>  Location: PIN_G19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[3]	=>  Location: PIN_R24,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[4]	=>  Location: PIN_H14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[5]	=>  Location: PIN_AF13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[6]	=>  Location: PIN_Y13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[7]	=>  Location: PIN_E14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[8]	=>  Location: PIN_A12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[9]	=>  Location: PIN_AF14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[10]	=>  Location: PIN_AC12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[11]	=>  Location: PIN_AE14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[12]	=>  Location: PIN_H19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[13]	=>  Location: PIN_AG18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[14]	=>  Location: PIN_G14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[15]	=>  Location: PIN_AD14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[16]	=>  Location: PIN_W22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[17]	=>  Location: PIN_AA12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[18]	=>  Location: PIN_F14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[19]	=>  Location: PIN_B11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[20]	=>  Location: PIN_A11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[21]	=>  Location: PIN_R28,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[22]	=>  Location: PIN_J14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[23]	=>  Location: PIN_AB13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[24]	=>  Location: PIN_N21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[25]	=>  Location: PIN_G22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[26]	=>  Location: PIN_F11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[27]	=>  Location: PIN_J13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[28]	=>  Location: PIN_F15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[29]	=>  Location: PIN_J16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[30]	=>  Location: PIN_AH18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[31]	=>  Location: PIN_AG17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tms	=>  Location: PIN_P8,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tck	=>  Location: PIN_P5,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdi	=>  Location: PIN_P7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdo	=>  Location: PIN_P6,	 I/O Standard: 2.5 V,	 Current Strength: Default


wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ;
wire \CPU|DP|dpif.halt~q ;
wire \CPU|DP|RU|reg_WEN~q ;
wire \CPU|DP|RU|reg_REN~q ;
wire \ramaddr~0_combout ;
wire \ramaddr~1_combout ;
wire \ramaddr~2_combout ;
wire \ramaddr~3_combout ;
wire \ramaddr~4_combout ;
wire \ramaddr~5_combout ;
wire \ramaddr~6_combout ;
wire \ramaddr~7_combout ;
wire \ramaddr~8_combout ;
wire \ramaddr~9_combout ;
wire \ramaddr~10_combout ;
wire \ramaddr~11_combout ;
wire \ramaddr~12_combout ;
wire \ramaddr~13_combout ;
wire \ramaddr~14_combout ;
wire \ramaddr~15_combout ;
wire \ramaddr~16_combout ;
wire \ramaddr~17_combout ;
wire \ramaddr~18_combout ;
wire \ramaddr~19_combout ;
wire \ramaddr~20_combout ;
wire \ramaddr~21_combout ;
wire \ramaddr~22_combout ;
wire \ramaddr~23_combout ;
wire \ramaddr~24_combout ;
wire \ramaddr~25_combout ;
wire \ramaddr~26_combout ;
wire \ramaddr~27_combout ;
wire \ramaddr~28_combout ;
wire \ramaddr~29_combout ;
wire \ramaddr~30_combout ;
wire \ramaddr~31_combout ;
wire \ramaddr~32_combout ;
wire \ramaddr~33_combout ;
wire \ramaddr~34_combout ;
wire \ramaddr~35_combout ;
wire \ramaddr~36_combout ;
wire \ramaddr~37_combout ;
wire \ramaddr~38_combout ;
wire \ramaddr~39_combout ;
wire \ramaddr~40_combout ;
wire \ramaddr~41_combout ;
wire \ramaddr~42_combout ;
wire \ramaddr~43_combout ;
wire \ramaddr~44_combout ;
wire \ramaddr~45_combout ;
wire \ramaddr~46_combout ;
wire \ramaddr~47_combout ;
wire \ramaddr~48_combout ;
wire \ramaddr~49_combout ;
wire \ramaddr~50_combout ;
wire \ramaddr~51_combout ;
wire \ramaddr~52_combout ;
wire \ramaddr~53_combout ;
wire \ramaddr~54_combout ;
wire \ramaddr~55_combout ;
wire \ramaddr~56_combout ;
wire \ramaddr~57_combout ;
wire \ramaddr~58_combout ;
wire \ramaddr~59_combout ;
wire \ramaddr~60_combout ;
wire \ramaddr~61_combout ;
wire \ramaddr~62_combout ;
wire \ramaddr~63_combout ;
wire \ramWEN~0_combout ;
wire \ramREN~0_combout ;
wire \RAM|always1~0_combout ;
wire \RAM|ramif.ramload[0]~0_combout ;
wire \RAM|ramif.ramload[1]~1_combout ;
wire \RAM|ramif.ramload[2]~2_combout ;
wire \RAM|ramif.ramload[3]~3_combout ;
wire \RAM|ramif.ramload[4]~4_combout ;
wire \RAM|ramif.ramload[5]~5_combout ;
wire \RAM|ramif.ramload[6]~6_combout ;
wire \RAM|ramif.ramload[7]~7_combout ;
wire \RAM|ramif.ramload[8]~8_combout ;
wire \RAM|ramif.ramload[9]~9_combout ;
wire \RAM|ramif.ramload[10]~10_combout ;
wire \RAM|ramif.ramload[11]~11_combout ;
wire \RAM|ramif.ramload[12]~12_combout ;
wire \RAM|ramif.ramload[13]~13_combout ;
wire \RAM|ramif.ramload[14]~14_combout ;
wire \RAM|ramif.ramload[15]~15_combout ;
wire \RAM|ramif.ramload[16]~17_combout ;
wire \RAM|ramif.ramload[17]~19_combout ;
wire \RAM|ramif.ramload[18]~20_combout ;
wire \RAM|ramif.ramload[19]~21_combout ;
wire \RAM|ramif.ramload[20]~22_combout ;
wire \RAM|ramif.ramload[21]~23_combout ;
wire \RAM|ramif.ramload[22]~24_combout ;
wire \RAM|ramif.ramload[23]~25_combout ;
wire \RAM|ramif.ramload[24]~26_combout ;
wire \RAM|ramif.ramload[25]~27_combout ;
wire \RAM|ramif.ramload[26]~28_combout ;
wire \RAM|ramif.ramload[27]~29_combout ;
wire \RAM|ramif.ramload[28]~30_combout ;
wire \RAM|ramif.ramload[29]~31_combout ;
wire \RAM|ramif.ramload[30]~32_combout ;
wire \RAM|ramif.ramload[31]~33_combout ;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ;
wire \CPUCLK~q ;
wire \CPU|DP|RF|Mux63~9_combout ;
wire \CPU|DP|RF|Mux63~23_combout ;
wire \CPU|CM|dcif.imemload[20]~10_combout ;
wire \ramstore~0_combout ;
wire \ramstore~1_combout ;
wire \CPU|DP|RF|Mux32~9_combout ;
wire \CPU|DP|RF|Mux32~19_combout ;
wire \CPU|DP|RF|Mux33~9_combout ;
wire \CPU|DP|RF|Mux33~19_combout ;
wire \CPU|DP|RF|Mux34~9_combout ;
wire \CPU|DP|RF|Mux34~19_combout ;
wire \CPU|DP|RF|Mux35~9_combout ;
wire \CPU|DP|RF|Mux35~19_combout ;
wire \CPU|DP|RF|Mux36~9_combout ;
wire \CPU|DP|RF|Mux36~19_combout ;
wire \CPU|DP|RF|Mux37~9_combout ;
wire \CPU|DP|RF|Mux37~19_combout ;
wire \CPU|DP|RF|Mux38~9_combout ;
wire \CPU|DP|RF|Mux38~19_combout ;
wire \CPU|DP|RF|Mux39~9_combout ;
wire \CPU|DP|RF|Mux39~19_combout ;
wire \CPU|DP|RF|Mux40~9_combout ;
wire \CPU|DP|RF|Mux40~19_combout ;
wire \CPU|DP|RF|Mux41~9_combout ;
wire \CPU|DP|RF|Mux41~19_combout ;
wire \CPU|DP|RF|Mux42~9_combout ;
wire \CPU|DP|RF|Mux42~19_combout ;
wire \CPU|DP|RF|Mux43~9_combout ;
wire \CPU|DP|RF|Mux43~19_combout ;
wire \CPU|DP|RF|Mux44~9_combout ;
wire \CPU|DP|RF|Mux44~19_combout ;
wire \CPU|DP|RF|Mux45~9_combout ;
wire \CPU|DP|RF|Mux45~19_combout ;
wire \CPU|DP|RF|Mux46~9_combout ;
wire \CPU|DP|RF|Mux46~19_combout ;
wire \CPU|DP|RF|Mux47~9_combout ;
wire \CPU|DP|RF|Mux47~19_combout ;
wire \CPU|DP|RF|Mux48~9_combout ;
wire \CPU|DP|RF|Mux48~19_combout ;
wire \CPU|DP|RF|Mux49~9_combout ;
wire \CPU|DP|RF|Mux49~19_combout ;
wire \CPU|DP|RF|Mux50~9_combout ;
wire \CPU|DP|RF|Mux50~19_combout ;
wire \CPU|DP|RF|Mux51~9_combout ;
wire \CPU|DP|RF|Mux51~19_combout ;
wire \CPU|DP|RF|Mux52~9_combout ;
wire \CPU|DP|RF|Mux52~19_combout ;
wire \CPU|DP|RF|Mux53~9_combout ;
wire \CPU|DP|RF|Mux53~19_combout ;
wire \CPU|DP|RF|Mux54~9_combout ;
wire \CPU|DP|RF|Mux54~19_combout ;
wire \CPU|DP|RF|Mux55~9_combout ;
wire \CPU|DP|RF|Mux55~19_combout ;
wire \CPU|DP|RF|Mux56~9_combout ;
wire \CPU|DP|RF|Mux56~19_combout ;
wire \CPU|DP|RF|Mux57~9_combout ;
wire \CPU|DP|RF|Mux57~19_combout ;
wire \CPU|DP|RF|Mux58~9_combout ;
wire \CPU|DP|RF|Mux58~19_combout ;
wire \CPU|DP|RF|Mux59~9_combout ;
wire \CPU|DP|RF|Mux59~19_combout ;
wire \CPU|DP|RF|Mux60~9_combout ;
wire \CPU|DP|RF|Mux60~19_combout ;
wire \CPU|DP|RF|Mux61~9_combout ;
wire \CPU|DP|RF|Mux61~19_combout ;
wire \CPU|DP|RF|Mux62~9_combout ;
wire \CPU|DP|RF|Mux62~21_combout ;
wire \ramstore~2_combout ;
wire \ramstore~3_combout ;
wire \ramstore~4_combout ;
wire \ramstore~5_combout ;
wire \ramstore~6_combout ;
wire \ramstore~7_combout ;
wire \ramstore~8_combout ;
wire \ramstore~9_combout ;
wire \ramstore~10_combout ;
wire \ramstore~11_combout ;
wire \ramstore~12_combout ;
wire \ramstore~13_combout ;
wire \ramstore~14_combout ;
wire \ramstore~15_combout ;
wire \ramstore~16_combout ;
wire \ramstore~17_combout ;
wire \ramstore~18_combout ;
wire \ramstore~19_combout ;
wire \ramstore~20_combout ;
wire \ramstore~21_combout ;
wire \ramstore~22_combout ;
wire \ramstore~23_combout ;
wire \ramstore~24_combout ;
wire \ramstore~25_combout ;
wire \ramstore~26_combout ;
wire \ramstore~27_combout ;
wire \ramstore~28_combout ;
wire \ramstore~29_combout ;
wire \ramstore~30_combout ;
wire \ramstore~31_combout ;
wire \ramstore~32_combout ;
wire \ramstore~33_combout ;
wire \ramstore~34_combout ;
wire \ramstore~35_combout ;
wire \ramstore~36_combout ;
wire \ramstore~37_combout ;
wire \ramstore~38_combout ;
wire \ramstore~39_combout ;
wire \ramstore~40_combout ;
wire \ramstore~41_combout ;
wire \ramstore~42_combout ;
wire \ramstore~43_combout ;
wire \ramstore~44_combout ;
wire \ramstore~45_combout ;
wire \ramstore~46_combout ;
wire \ramstore~47_combout ;
wire \ramstore~48_combout ;
wire \ramstore~49_combout ;
wire \ramstore~50_combout ;
wire \ramstore~51_combout ;
wire \ramstore~52_combout ;
wire \ramstore~53_combout ;
wire \ramstore~54_combout ;
wire \ramstore~55_combout ;
wire \ramstore~56_combout ;
wire \ramstore~57_combout ;
wire \ramstore~58_combout ;
wire \ramstore~59_combout ;
wire \ramstore~60_combout ;
wire \ramstore~61_combout ;
wire \ramstore~62_combout ;
wire \ramstore~63_combout ;
wire \Equal0~0_combout ;
wire \CPUCLK~0_combout ;
wire \count[3]~0_combout ;
wire \count[2]~1_combout ;
wire \count[1]~2_combout ;
wire \count~3_combout ;
wire \ramaddr~29_wirecell_combout ;
wire \altera_internal_jtag~TCKUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ;
wire \syif.tbCTRL~input_o ;
wire \syif.addr[1]~input_o ;
wire \syif.addr[0]~input_o ;
wire \syif.addr[3]~input_o ;
wire \syif.addr[2]~input_o ;
wire \syif.addr[5]~input_o ;
wire \syif.addr[4]~input_o ;
wire \syif.addr[7]~input_o ;
wire \syif.addr[6]~input_o ;
wire \syif.addr[9]~input_o ;
wire \syif.addr[8]~input_o ;
wire \syif.addr[11]~input_o ;
wire \syif.addr[10]~input_o ;
wire \syif.addr[13]~input_o ;
wire \syif.addr[12]~input_o ;
wire \syif.addr[15]~input_o ;
wire \syif.addr[14]~input_o ;
wire \syif.addr[17]~input_o ;
wire \syif.addr[16]~input_o ;
wire \syif.addr[19]~input_o ;
wire \syif.addr[18]~input_o ;
wire \syif.addr[21]~input_o ;
wire \syif.addr[20]~input_o ;
wire \syif.addr[23]~input_o ;
wire \syif.addr[22]~input_o ;
wire \syif.addr[25]~input_o ;
wire \syif.addr[24]~input_o ;
wire \syif.addr[27]~input_o ;
wire \syif.addr[26]~input_o ;
wire \syif.addr[29]~input_o ;
wire \syif.addr[28]~input_o ;
wire \syif.addr[31]~input_o ;
wire \syif.addr[30]~input_o ;
wire \syif.WEN~input_o ;
wire \syif.REN~input_o ;
wire \nRST~input_o ;
wire \CLK~input_o ;
wire \syif.store[0]~input_o ;
wire \syif.store[1]~input_o ;
wire \syif.store[2]~input_o ;
wire \syif.store[3]~input_o ;
wire \syif.store[4]~input_o ;
wire \syif.store[5]~input_o ;
wire \syif.store[6]~input_o ;
wire \syif.store[7]~input_o ;
wire \syif.store[8]~input_o ;
wire \syif.store[9]~input_o ;
wire \syif.store[10]~input_o ;
wire \syif.store[11]~input_o ;
wire \syif.store[12]~input_o ;
wire \syif.store[13]~input_o ;
wire \syif.store[14]~input_o ;
wire \syif.store[15]~input_o ;
wire \syif.store[16]~input_o ;
wire \syif.store[17]~input_o ;
wire \syif.store[18]~input_o ;
wire \syif.store[19]~input_o ;
wire \syif.store[20]~input_o ;
wire \syif.store[21]~input_o ;
wire \syif.store[22]~input_o ;
wire \syif.store[23]~input_o ;
wire \syif.store[24]~input_o ;
wire \syif.store[25]~input_o ;
wire \syif.store[26]~input_o ;
wire \syif.store[27]~input_o ;
wire \syif.store[28]~input_o ;
wire \syif.store[29]~input_o ;
wire \syif.store[30]~input_o ;
wire \syif.store[31]~input_o ;
wire \altera_internal_jtag~TCKUTAPclkctrl_outclk ;
wire \CPUCLK~clkctrl_outclk ;
wire \nRST~inputclkctrl_outclk ;
wire \CLK~inputclkctrl_outclk ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~10 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13_combout ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ;
wire \~QIC_CREATED_GND~I_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ;
wire \altera_internal_jtag~TDO ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg ;
wire [9:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg ;
wire [5:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt ;
wire [15:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR ;
wire [3:0] count;
wire [31:0] \CPU|DP|PCU|PC ;
wire [31:0] \CPU|CM|daddr ;
wire [3:0] \RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg ;


ram RAM(
	.is_in_use_reg(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.ramaddr(\ramaddr~1_combout ),
	.ramaddr1(\ramaddr~3_combout ),
	.ramaddr2(\ramaddr~5_combout ),
	.ramaddr3(\ramaddr~7_combout ),
	.ramaddr4(\ramaddr~9_combout ),
	.ramaddr5(\ramaddr~11_combout ),
	.ramaddr6(\ramaddr~13_combout ),
	.ramaddr7(\ramaddr~15_combout ),
	.ramaddr8(\ramaddr~17_combout ),
	.ramaddr9(\ramaddr~19_combout ),
	.ramaddr10(\ramaddr~21_combout ),
	.ramaddr11(\ramaddr~23_combout ),
	.ramaddr12(\ramaddr~25_combout ),
	.ramaddr13(\ramaddr~27_combout ),
	.ramaddr14(\ramaddr~29_combout ),
	.ramaddr15(\ramaddr~31_combout ),
	.\ramif.ramaddr ({\ramaddr~61_combout ,gnd,\ramaddr~57_combout ,gnd,\ramaddr~53_combout ,gnd,gnd,gnd,\ramaddr~45_combout ,gnd,\ramaddr~41_combout ,gnd,\ramaddr~37_combout ,gnd,\ramaddr~33_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.ramaddr16(\ramaddr~35_combout ),
	.ramaddr17(\ramaddr~39_combout ),
	.ramaddr18(\ramaddr~43_combout ),
	.ramaddr19(\ramaddr~47_combout ),
	.ramaddr20(\ramaddr~49_combout ),
	.ramaddr21(\ramaddr~51_combout ),
	.ramaddr22(\ramaddr~55_combout ),
	.ramaddr23(\ramaddr~59_combout ),
	.ramaddr24(\ramaddr~63_combout ),
	.\ramif.ramWEN (\ramWEN~0_combout ),
	.\ramif.ramREN (\ramREN~0_combout ),
	.always1(\RAM|always1~0_combout ),
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~1_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~2_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~3_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~4_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~5_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~6_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~7_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~8_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~9_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~10_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~11_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~12_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~13_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~14_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~15_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~17_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~19_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~20_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~21_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~22_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~23_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~24_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~25_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~26_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~27_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~28_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~29_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~30_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~31_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~32_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~33_combout ),
	.ir_loaded_address_reg_0(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.ir_loaded_address_reg_1(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.ir_loaded_address_reg_2(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.ir_loaded_address_reg_3(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.tdo(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.ramstore(\ramstore~1_combout ),
	.ramstore1(\ramstore~3_combout ),
	.ramstore2(\ramstore~5_combout ),
	.ramstore3(\ramstore~7_combout ),
	.ramstore4(\ramstore~9_combout ),
	.ramstore5(\ramstore~11_combout ),
	.ramstore6(\ramstore~13_combout ),
	.ramstore7(\ramstore~15_combout ),
	.ramstore8(\ramstore~17_combout ),
	.ramstore9(\ramstore~19_combout ),
	.ramstore10(\ramstore~21_combout ),
	.ramstore11(\ramstore~23_combout ),
	.ramstore12(\ramstore~25_combout ),
	.ramstore13(\ramstore~27_combout ),
	.ramstore14(\ramstore~29_combout ),
	.ramstore15(\ramstore~31_combout ),
	.ramstore16(\ramstore~33_combout ),
	.ramstore17(\ramstore~35_combout ),
	.ramstore18(\ramstore~37_combout ),
	.ramstore19(\ramstore~39_combout ),
	.ramstore20(\ramstore~41_combout ),
	.ramstore21(\ramstore~43_combout ),
	.ramstore22(\ramstore~45_combout ),
	.ramstore23(\ramstore~47_combout ),
	.ramstore24(\ramstore~49_combout ),
	.ramstore25(\ramstore~51_combout ),
	.ramstore26(\ramstore~53_combout ),
	.ramstore27(\ramstore~55_combout ),
	.ramstore28(\ramstore~57_combout ),
	.ramstore29(\ramstore~59_combout ),
	.ramstore30(\ramstore~61_combout ),
	.ramstore31(\ramstore~63_combout ),
	.ramaddr25(\ramaddr~29_wirecell_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.irf_reg_0_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.irf_reg_1_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.irf_reg_2_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.irf_reg_3_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.irf_reg_4_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.node_ena_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.clr_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.virtual_ir_scan_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.state_5(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.state_8(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.nRST(\nRST~input_o ),
	.altera_internal_jtag1(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.nRST1(\nRST~inputclkctrl_outclk ),
	.CLK(\CLK~inputclkctrl_outclk ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

singlecycle CPU(
	.PC_29(\CPU|DP|PCU|PC [29]),
	.PC_28(\CPU|DP|PCU|PC [28]),
	.PC_31(\CPU|DP|PCU|PC [31]),
	.PC_30(\CPU|DP|PCU|PC [30]),
	.dpifhalt(\CPU|DP|dpif.halt~q ),
	.PC_1(\CPU|DP|PCU|PC [1]),
	.daddr_1(\CPU|CM|daddr [1]),
	.reg_WEN(\CPU|DP|RU|reg_WEN~q ),
	.reg_REN(\CPU|DP|RU|reg_REN~q ),
	.PC_0(\CPU|DP|PCU|PC [0]),
	.daddr_0(\CPU|CM|daddr [0]),
	.daddr_3(\CPU|CM|daddr [3]),
	.PC_3(\CPU|DP|PCU|PC [3]),
	.daddr_2(\CPU|CM|daddr [2]),
	.PC_2(\CPU|DP|PCU|PC [2]),
	.daddr_5(\CPU|CM|daddr [5]),
	.PC_5(\CPU|DP|PCU|PC [5]),
	.PC_4(\CPU|DP|PCU|PC [4]),
	.daddr_4(\CPU|CM|daddr [4]),
	.PC_7(\CPU|DP|PCU|PC [7]),
	.daddr_7(\CPU|CM|daddr [7]),
	.daddr_6(\CPU|CM|daddr [6]),
	.PC_6(\CPU|DP|PCU|PC [6]),
	.daddr_9(\CPU|CM|daddr [9]),
	.PC_9(\CPU|DP|PCU|PC [9]),
	.daddr_8(\CPU|CM|daddr [8]),
	.PC_8(\CPU|DP|PCU|PC [8]),
	.daddr_11(\CPU|CM|daddr [11]),
	.PC_11(\CPU|DP|PCU|PC [11]),
	.daddr_10(\CPU|CM|daddr [10]),
	.PC_10(\CPU|DP|PCU|PC [10]),
	.PC_13(\CPU|DP|PCU|PC [13]),
	.daddr_13(\CPU|CM|daddr [13]),
	.daddr_12(\CPU|CM|daddr [12]),
	.PC_12(\CPU|DP|PCU|PC [12]),
	.daddr_15(\CPU|CM|daddr [15]),
	.PC_15(\CPU|DP|PCU|PC [15]),
	.daddr_14(\CPU|CM|daddr [14]),
	.PC_14(\CPU|DP|PCU|PC [14]),
	.daddr_17(\CPU|CM|daddr [17]),
	.PC_17(\CPU|DP|PCU|PC [17]),
	.PC_16(\CPU|DP|PCU|PC [16]),
	.daddr_16(\CPU|CM|daddr [16]),
	.daddr_19(\CPU|CM|daddr [19]),
	.PC_19(\CPU|DP|PCU|PC [19]),
	.daddr_18(\CPU|CM|daddr [18]),
	.PC_18(\CPU|DP|PCU|PC [18]),
	.PC_21(\CPU|DP|PCU|PC [21]),
	.daddr_21(\CPU|CM|daddr [21]),
	.daddr_20(\CPU|CM|daddr [20]),
	.PC_20(\CPU|DP|PCU|PC [20]),
	.daddr_23(\CPU|CM|daddr [23]),
	.PC_23(\CPU|DP|PCU|PC [23]),
	.daddr_22(\CPU|CM|daddr [22]),
	.PC_22(\CPU|DP|PCU|PC [22]),
	.daddr_25(\CPU|CM|daddr [25]),
	.PC_25(\CPU|DP|PCU|PC [25]),
	.daddr_24(\CPU|CM|daddr [24]),
	.PC_24(\CPU|DP|PCU|PC [24]),
	.PC_27(\CPU|DP|PCU|PC [27]),
	.daddr_27(\CPU|CM|daddr [27]),
	.daddr_26(\CPU|CM|daddr [26]),
	.PC_26(\CPU|DP|PCU|PC [26]),
	.daddr_29(\CPU|CM|daddr [29]),
	.daddr_28(\CPU|CM|daddr [28]),
	.daddr_31(\CPU|CM|daddr [31]),
	.daddr_30(\CPU|CM|daddr [30]),
	.always1(\RAM|always1~0_combout ),
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~1_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~2_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~3_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~4_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~5_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~6_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~7_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~8_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~9_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~10_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~11_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~12_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~13_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~14_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~15_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~17_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~19_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~20_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~21_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~22_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~23_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~24_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~25_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~26_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~27_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~28_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~29_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~30_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~31_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~32_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~33_combout ),
	.Mux63(\CPU|DP|RF|Mux63~9_combout ),
	.Mux631(\CPU|DP|RF|Mux63~23_combout ),
	.dcifimemload_20(\CPU|CM|dcif.imemload[20]~10_combout ),
	.Mux32(\CPU|DP|RF|Mux32~9_combout ),
	.Mux321(\CPU|DP|RF|Mux32~19_combout ),
	.Mux33(\CPU|DP|RF|Mux33~9_combout ),
	.Mux331(\CPU|DP|RF|Mux33~19_combout ),
	.Mux34(\CPU|DP|RF|Mux34~9_combout ),
	.Mux341(\CPU|DP|RF|Mux34~19_combout ),
	.Mux35(\CPU|DP|RF|Mux35~9_combout ),
	.Mux351(\CPU|DP|RF|Mux35~19_combout ),
	.Mux36(\CPU|DP|RF|Mux36~9_combout ),
	.Mux361(\CPU|DP|RF|Mux36~19_combout ),
	.Mux37(\CPU|DP|RF|Mux37~9_combout ),
	.Mux371(\CPU|DP|RF|Mux37~19_combout ),
	.Mux38(\CPU|DP|RF|Mux38~9_combout ),
	.Mux381(\CPU|DP|RF|Mux38~19_combout ),
	.Mux39(\CPU|DP|RF|Mux39~9_combout ),
	.Mux391(\CPU|DP|RF|Mux39~19_combout ),
	.Mux40(\CPU|DP|RF|Mux40~9_combout ),
	.Mux401(\CPU|DP|RF|Mux40~19_combout ),
	.Mux41(\CPU|DP|RF|Mux41~9_combout ),
	.Mux411(\CPU|DP|RF|Mux41~19_combout ),
	.Mux42(\CPU|DP|RF|Mux42~9_combout ),
	.Mux421(\CPU|DP|RF|Mux42~19_combout ),
	.Mux43(\CPU|DP|RF|Mux43~9_combout ),
	.Mux431(\CPU|DP|RF|Mux43~19_combout ),
	.Mux44(\CPU|DP|RF|Mux44~9_combout ),
	.Mux441(\CPU|DP|RF|Mux44~19_combout ),
	.Mux45(\CPU|DP|RF|Mux45~9_combout ),
	.Mux451(\CPU|DP|RF|Mux45~19_combout ),
	.Mux46(\CPU|DP|RF|Mux46~9_combout ),
	.Mux461(\CPU|DP|RF|Mux46~19_combout ),
	.Mux47(\CPU|DP|RF|Mux47~9_combout ),
	.Mux471(\CPU|DP|RF|Mux47~19_combout ),
	.Mux48(\CPU|DP|RF|Mux48~9_combout ),
	.Mux481(\CPU|DP|RF|Mux48~19_combout ),
	.Mux49(\CPU|DP|RF|Mux49~9_combout ),
	.Mux491(\CPU|DP|RF|Mux49~19_combout ),
	.Mux50(\CPU|DP|RF|Mux50~9_combout ),
	.Mux501(\CPU|DP|RF|Mux50~19_combout ),
	.Mux51(\CPU|DP|RF|Mux51~9_combout ),
	.Mux511(\CPU|DP|RF|Mux51~19_combout ),
	.Mux52(\CPU|DP|RF|Mux52~9_combout ),
	.Mux521(\CPU|DP|RF|Mux52~19_combout ),
	.Mux53(\CPU|DP|RF|Mux53~9_combout ),
	.Mux531(\CPU|DP|RF|Mux53~19_combout ),
	.Mux54(\CPU|DP|RF|Mux54~9_combout ),
	.Mux541(\CPU|DP|RF|Mux54~19_combout ),
	.Mux55(\CPU|DP|RF|Mux55~9_combout ),
	.Mux551(\CPU|DP|RF|Mux55~19_combout ),
	.Mux56(\CPU|DP|RF|Mux56~9_combout ),
	.Mux561(\CPU|DP|RF|Mux56~19_combout ),
	.Mux57(\CPU|DP|RF|Mux57~9_combout ),
	.Mux571(\CPU|DP|RF|Mux57~19_combout ),
	.Mux58(\CPU|DP|RF|Mux58~9_combout ),
	.Mux581(\CPU|DP|RF|Mux58~19_combout ),
	.Mux59(\CPU|DP|RF|Mux59~9_combout ),
	.Mux591(\CPU|DP|RF|Mux59~19_combout ),
	.Mux60(\CPU|DP|RF|Mux60~9_combout ),
	.Mux601(\CPU|DP|RF|Mux60~19_combout ),
	.Mux61(\CPU|DP|RF|Mux61~9_combout ),
	.Mux611(\CPU|DP|RF|Mux61~19_combout ),
	.Mux62(\CPU|DP|RF|Mux62~9_combout ),
	.Mux621(\CPU|DP|RF|Mux62~21_combout ),
	.nRST(\nRST~input_o ),
	.CLK(\CPUCLK~clkctrl_outclk ),
	.nRST1(\nRST~inputclkctrl_outclk ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X60_Y33_N30
cycloneive_lcell_comb \ramaddr~0 (
// Equation(s):
// \ramaddr~0_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[1]~input_o )) # (!\syif.tbCTRL~input_o  & (((!reg_REN1 & !reg_WEN1))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[1]~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramaddr~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~0 .lut_mask = 16'h888D;
defparam \ramaddr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N12
cycloneive_lcell_comb \ramaddr~1 (
// Equation(s):
// \ramaddr~1_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~0_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~0_combout  & ((PC_1))) # (!\ramaddr~0_combout  & (daddr_1))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [1]),
	.datac(\ramaddr~0_combout ),
	.datad(\CPU|DP|PCU|PC [1]),
	.cin(gnd),
	.combout(\ramaddr~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~1 .lut_mask = 16'hF4A4;
defparam \ramaddr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N28
cycloneive_lcell_comb \ramaddr~2 (
// Equation(s):
// \ramaddr~2_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[0]~input_o )) # (!\syif.tbCTRL~input_o  & (((!reg_REN1 & !reg_WEN1))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[0]~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramaddr~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~2 .lut_mask = 16'h888D;
defparam \ramaddr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N6
cycloneive_lcell_comb \ramaddr~3 (
// Equation(s):
// \ramaddr~3_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~2_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~2_combout  & (PC_0)) # (!\ramaddr~2_combout  & ((daddr_0)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|PCU|PC [0]),
	.datac(\CPU|CM|daddr [0]),
	.datad(\ramaddr~2_combout ),
	.cin(gnd),
	.combout(\ramaddr~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~3 .lut_mask = 16'hEE50;
defparam \ramaddr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N2
cycloneive_lcell_comb \ramaddr~4 (
// Equation(s):
// \ramaddr~4_combout  = (reg_WEN1 & (daddr_3)) # (!reg_WEN1 & ((reg_REN1 & (daddr_3)) # (!reg_REN1 & ((PC_3)))))

	.dataa(\CPU|CM|daddr [3]),
	.datab(\CPU|DP|PCU|PC [3]),
	.datac(\CPU|DP|RU|reg_WEN~q ),
	.datad(\CPU|DP|RU|reg_REN~q ),
	.cin(gnd),
	.combout(\ramaddr~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~4 .lut_mask = 16'hAAAC;
defparam \ramaddr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N0
cycloneive_lcell_comb \ramaddr~5 (
// Equation(s):
// \ramaddr~5_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[3]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~4_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[3]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~4_combout ),
	.cin(gnd),
	.combout(\ramaddr~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~5 .lut_mask = 16'hDD88;
defparam \ramaddr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N20
cycloneive_lcell_comb \ramaddr~6 (
// Equation(s):
// \ramaddr~6_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[2]~input_o )) # (!\syif.tbCTRL~input_o  & (((reg_WEN1) # (reg_REN1))))

	.dataa(\syif.addr[2]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RU|reg_WEN~q ),
	.datad(\CPU|DP|RU|reg_REN~q ),
	.cin(gnd),
	.combout(\ramaddr~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~6 .lut_mask = 16'hBBB8;
defparam \ramaddr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N10
cycloneive_lcell_comb \ramaddr~7 (
// Equation(s):
// \ramaddr~7_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~6_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~6_combout  & (daddr_2)) # (!\ramaddr~6_combout  & ((PC_2)))))

	.dataa(\CPU|CM|daddr [2]),
	.datab(\CPU|DP|PCU|PC [2]),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~6_combout ),
	.cin(gnd),
	.combout(\ramaddr~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~7 .lut_mask = 16'hFA0C;
defparam \ramaddr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N8
cycloneive_lcell_comb \ramaddr~8 (
// Equation(s):
// \ramaddr~8_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[5]~input_o )))) # (!\syif.tbCTRL~input_o  & ((reg_WEN1) # ((reg_REN1))))

	.dataa(\CPU|DP|RU|reg_WEN~q ),
	.datab(\syif.addr[5]~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramaddr~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~8 .lut_mask = 16'hCCFA;
defparam \ramaddr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N22
cycloneive_lcell_comb \ramaddr~9 (
// Equation(s):
// \ramaddr~9_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~8_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~8_combout  & ((daddr_5))) # (!\ramaddr~8_combout  & (PC_5))))

	.dataa(\CPU|DP|PCU|PC [5]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramaddr~8_combout ),
	.datad(\CPU|CM|daddr [5]),
	.cin(gnd),
	.combout(\ramaddr~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~9 .lut_mask = 16'hF2C2;
defparam \ramaddr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N26
cycloneive_lcell_comb \ramaddr~10 (
// Equation(s):
// \ramaddr~10_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[4]~input_o )))) # (!\syif.tbCTRL~input_o  & (!reg_WEN1 & ((!reg_REN1))))

	.dataa(\CPU|DP|RU|reg_WEN~q ),
	.datab(\syif.addr[4]~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramaddr~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~10 .lut_mask = 16'hCC05;
defparam \ramaddr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N24
cycloneive_lcell_comb \ramaddr~11 (
// Equation(s):
// \ramaddr~11_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~10_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~10_combout  & (PC_4)) # (!\ramaddr~10_combout  & ((daddr_4)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|PCU|PC [4]),
	.datac(\ramaddr~10_combout ),
	.datad(\CPU|CM|daddr [4]),
	.cin(gnd),
	.combout(\ramaddr~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~11 .lut_mask = 16'hE5E0;
defparam \ramaddr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N18
cycloneive_lcell_comb \ramaddr~12 (
// Equation(s):
// \ramaddr~12_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[7]~input_o )) # (!\syif.tbCTRL~input_o  & (((!reg_WEN1 & !reg_REN1))))

	.dataa(\syif.addr[7]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RU|reg_WEN~q ),
	.datad(\CPU|DP|RU|reg_REN~q ),
	.cin(gnd),
	.combout(\ramaddr~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~12 .lut_mask = 16'h888B;
defparam \ramaddr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N16
cycloneive_lcell_comb \ramaddr~13 (
// Equation(s):
// \ramaddr~13_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~12_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~12_combout  & (PC_7)) # (!\ramaddr~12_combout  & ((daddr_7)))))

	.dataa(\CPU|DP|PCU|PC [7]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|CM|daddr [7]),
	.datad(\ramaddr~12_combout ),
	.cin(gnd),
	.combout(\ramaddr~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~13 .lut_mask = 16'hEE30;
defparam \ramaddr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N6
cycloneive_lcell_comb \ramaddr~14 (
// Equation(s):
// \ramaddr~14_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[6]~input_o )) # (!\syif.tbCTRL~input_o  & (((reg_WEN1) # (reg_REN1))))

	.dataa(\syif.addr[6]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RU|reg_WEN~q ),
	.datad(\CPU|DP|RU|reg_REN~q ),
	.cin(gnd),
	.combout(\ramaddr~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~14 .lut_mask = 16'hBBB8;
defparam \ramaddr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N20
cycloneive_lcell_comb \ramaddr~15 (
// Equation(s):
// \ramaddr~15_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~14_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~14_combout  & (daddr_6)) # (!\ramaddr~14_combout  & ((PC_6)))))

	.dataa(\CPU|CM|daddr [6]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|PCU|PC [6]),
	.datad(\ramaddr~14_combout ),
	.cin(gnd),
	.combout(\ramaddr~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~15 .lut_mask = 16'hEE30;
defparam \ramaddr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N6
cycloneive_lcell_comb \ramaddr~16 (
// Equation(s):
// \ramaddr~16_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[9]~input_o )) # (!\syif.tbCTRL~input_o  & (((reg_REN1) # (reg_WEN1))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[9]~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramaddr~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~16 .lut_mask = 16'hDDD8;
defparam \ramaddr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N24
cycloneive_lcell_comb \ramaddr~17 (
// Equation(s):
// \ramaddr~17_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~16_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~16_combout  & (daddr_9)) # (!\ramaddr~16_combout  & ((PC_9)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [9]),
	.datac(\CPU|DP|PCU|PC [9]),
	.datad(\ramaddr~16_combout ),
	.cin(gnd),
	.combout(\ramaddr~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~17 .lut_mask = 16'hEE50;
defparam \ramaddr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N12
cycloneive_lcell_comb \ramaddr~18 (
// Equation(s):
// \ramaddr~18_combout  = (reg_REN1 & (((daddr_8)))) # (!reg_REN1 & ((reg_WEN1 & ((daddr_8))) # (!reg_WEN1 & (PC_8))))

	.dataa(\CPU|DP|PCU|PC [8]),
	.datab(\CPU|CM|daddr [8]),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramaddr~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~18 .lut_mask = 16'hCCCA;
defparam \ramaddr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N2
cycloneive_lcell_comb \ramaddr~19 (
// Equation(s):
// \ramaddr~19_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[8]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~18_combout )))

	.dataa(gnd),
	.datab(\syif.addr[8]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~18_combout ),
	.cin(gnd),
	.combout(\ramaddr~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~19 .lut_mask = 16'hCFC0;
defparam \ramaddr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N10
cycloneive_lcell_comb \ramaddr~20 (
// Equation(s):
// \ramaddr~20_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[11]~input_o )) # (!\syif.tbCTRL~input_o  & (((reg_REN1) # (reg_WEN1))))

	.dataa(\syif.addr[11]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramaddr~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~20 .lut_mask = 16'hBBB8;
defparam \ramaddr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N16
cycloneive_lcell_comb \ramaddr~21 (
// Equation(s):
// \ramaddr~21_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~20_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~20_combout  & (daddr_11)) # (!\ramaddr~20_combout  & ((PC_11)))))

	.dataa(\CPU|CM|daddr [11]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|PCU|PC [11]),
	.datad(\ramaddr~20_combout ),
	.cin(gnd),
	.combout(\ramaddr~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~21 .lut_mask = 16'hEE30;
defparam \ramaddr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N2
cycloneive_lcell_comb \ramaddr~22 (
// Equation(s):
// \ramaddr~22_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[10]~input_o )) # (!\syif.tbCTRL~input_o  & (((reg_REN1) # (reg_WEN1))))

	.dataa(\syif.addr[10]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramaddr~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~22 .lut_mask = 16'hBBB8;
defparam \ramaddr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N20
cycloneive_lcell_comb \ramaddr~23 (
// Equation(s):
// \ramaddr~23_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~22_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~22_combout  & ((daddr_10))) # (!\ramaddr~22_combout  & (PC_10))))

	.dataa(\CPU|DP|PCU|PC [10]),
	.datab(\CPU|CM|daddr [10]),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~22_combout ),
	.cin(gnd),
	.combout(\ramaddr~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~23 .lut_mask = 16'hFC0A;
defparam \ramaddr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N2
cycloneive_lcell_comb \ramaddr~24 (
// Equation(s):
// \ramaddr~24_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[13]~input_o )))) # (!\syif.tbCTRL~input_o  & (!reg_REN1 & (!reg_WEN1)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|RU|reg_REN~q ),
	.datac(\CPU|DP|RU|reg_WEN~q ),
	.datad(\syif.addr[13]~input_o ),
	.cin(gnd),
	.combout(\ramaddr~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~24 .lut_mask = 16'hAB01;
defparam \ramaddr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N24
cycloneive_lcell_comb \ramaddr~25 (
// Equation(s):
// \ramaddr~25_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~24_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~24_combout  & ((PC_13))) # (!\ramaddr~24_combout  & (daddr_13))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [13]),
	.datac(\CPU|DP|PCU|PC [13]),
	.datad(\ramaddr~24_combout ),
	.cin(gnd),
	.combout(\ramaddr~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~25 .lut_mask = 16'hFA44;
defparam \ramaddr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N16
cycloneive_lcell_comb \ramaddr~26 (
// Equation(s):
// \ramaddr~26_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[12]~input_o )))) # (!\syif.tbCTRL~input_o  & ((reg_REN1) # ((reg_WEN1))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|RU|reg_REN~q ),
	.datac(\CPU|DP|RU|reg_WEN~q ),
	.datad(\syif.addr[12]~input_o ),
	.cin(gnd),
	.combout(\ramaddr~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~26 .lut_mask = 16'hFE54;
defparam \ramaddr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N18
cycloneive_lcell_comb \ramaddr~27 (
// Equation(s):
// \ramaddr~27_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~26_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~26_combout  & (daddr_12)) # (!\ramaddr~26_combout  & ((PC_12)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [12]),
	.datac(\CPU|DP|PCU|PC [12]),
	.datad(\ramaddr~26_combout ),
	.cin(gnd),
	.combout(\ramaddr~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~27 .lut_mask = 16'hEE50;
defparam \ramaddr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N6
cycloneive_lcell_comb \ramaddr~28 (
// Equation(s):
// \ramaddr~28_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[15]~input_o )) # (!\syif.tbCTRL~input_o  & (((reg_REN1) # (reg_WEN1))))

	.dataa(\syif.addr[15]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramaddr~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~28 .lut_mask = 16'hBBB8;
defparam \ramaddr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N16
cycloneive_lcell_comb \ramaddr~29 (
// Equation(s):
// \ramaddr~29_combout  = (\syif.tbCTRL~input_o  & (((!\ramaddr~28_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~28_combout  & (!daddr_15)) # (!\ramaddr~28_combout  & ((!PC_15)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [15]),
	.datac(\CPU|DP|PCU|PC [15]),
	.datad(\ramaddr~28_combout ),
	.cin(gnd),
	.combout(\ramaddr~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29 .lut_mask = 16'h11AF;
defparam \ramaddr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N20
cycloneive_lcell_comb \ramaddr~30 (
// Equation(s):
// \ramaddr~30_combout  = (reg_WEN1 & (daddr_14)) # (!reg_WEN1 & ((reg_REN1 & (daddr_14)) # (!reg_REN1 & ((PC_14)))))

	.dataa(\CPU|DP|RU|reg_WEN~q ),
	.datab(\CPU|CM|daddr [14]),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|DP|PCU|PC [14]),
	.cin(gnd),
	.combout(\ramaddr~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~30 .lut_mask = 16'hCDC8;
defparam \ramaddr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N10
cycloneive_lcell_comb \ramaddr~31 (
// Equation(s):
// \ramaddr~31_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[14]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~30_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[14]~input_o ),
	.datad(\ramaddr~30_combout ),
	.cin(gnd),
	.combout(\ramaddr~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~31 .lut_mask = 16'hF3C0;
defparam \ramaddr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N2
cycloneive_lcell_comb \ramaddr~32 (
// Equation(s):
// \ramaddr~32_combout  = (reg_WEN1 & (((daddr_17)))) # (!reg_WEN1 & ((reg_REN1 & ((daddr_17))) # (!reg_REN1 & (PC_17))))

	.dataa(\CPU|DP|RU|reg_WEN~q ),
	.datab(\CPU|DP|PCU|PC [17]),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|CM|daddr [17]),
	.cin(gnd),
	.combout(\ramaddr~32_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~32 .lut_mask = 16'hFE04;
defparam \ramaddr~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N20
cycloneive_lcell_comb \ramaddr~33 (
// Equation(s):
// \ramaddr~33_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[17]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~32_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[17]~input_o ),
	.datad(\ramaddr~32_combout ),
	.cin(gnd),
	.combout(\ramaddr~33_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~33 .lut_mask = 16'hF3C0;
defparam \ramaddr~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N18
cycloneive_lcell_comb \ramaddr~34 (
// Equation(s):
// \ramaddr~34_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[16]~input_o )))) # (!\syif.tbCTRL~input_o  & (!reg_WEN1 & (!reg_REN1)))

	.dataa(\CPU|DP|RU|reg_WEN~q ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\syif.addr[16]~input_o ),
	.cin(gnd),
	.combout(\ramaddr~34_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~34 .lut_mask = 16'hCD01;
defparam \ramaddr~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N16
cycloneive_lcell_comb \ramaddr~35 (
// Equation(s):
// \ramaddr~35_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~34_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~34_combout  & (PC_16)) # (!\ramaddr~34_combout  & ((daddr_16)))))

	.dataa(\CPU|DP|PCU|PC [16]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|CM|daddr [16]),
	.datad(\ramaddr~34_combout ),
	.cin(gnd),
	.combout(\ramaddr~35_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~35 .lut_mask = 16'hEE30;
defparam \ramaddr~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N6
cycloneive_lcell_comb \ramaddr~36 (
// Equation(s):
// \ramaddr~36_combout  = (reg_REN1 & (((daddr_19)))) # (!reg_REN1 & ((reg_WEN1 & ((daddr_19))) # (!reg_WEN1 & (PC_19))))

	.dataa(\CPU|DP|RU|reg_REN~q ),
	.datab(\CPU|DP|PCU|PC [19]),
	.datac(\CPU|CM|daddr [19]),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramaddr~36_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~36 .lut_mask = 16'hF0E4;
defparam \ramaddr~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N12
cycloneive_lcell_comb \ramaddr~37 (
// Equation(s):
// \ramaddr~37_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[19]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~36_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[19]~input_o ),
	.datad(\ramaddr~36_combout ),
	.cin(gnd),
	.combout(\ramaddr~37_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~37 .lut_mask = 16'hF3C0;
defparam \ramaddr~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N0
cycloneive_lcell_comb \ramaddr~38 (
// Equation(s):
// \ramaddr~38_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[18]~input_o )))) # (!\syif.tbCTRL~input_o  & ((reg_WEN1) # ((reg_REN1))))

	.dataa(\CPU|DP|RU|reg_WEN~q ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\syif.addr[18]~input_o ),
	.cin(gnd),
	.combout(\ramaddr~38_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~38 .lut_mask = 16'hFE32;
defparam \ramaddr~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N30
cycloneive_lcell_comb \ramaddr~39 (
// Equation(s):
// \ramaddr~39_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~38_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~38_combout  & (daddr_18)) # (!\ramaddr~38_combout  & ((PC_18)))))

	.dataa(\CPU|CM|daddr [18]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|PCU|PC [18]),
	.datad(\ramaddr~38_combout ),
	.cin(gnd),
	.combout(\ramaddr~39_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~39 .lut_mask = 16'hEE30;
defparam \ramaddr~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N12
cycloneive_lcell_comb \ramaddr~40 (
// Equation(s):
// \ramaddr~40_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[21]~input_o )) # (!\syif.tbCTRL~input_o  & (((!reg_WEN1 & !reg_REN1))))

	.dataa(\syif.addr[21]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RU|reg_WEN~q ),
	.datad(\CPU|DP|RU|reg_REN~q ),
	.cin(gnd),
	.combout(\ramaddr~40_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~40 .lut_mask = 16'h888B;
defparam \ramaddr~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N14
cycloneive_lcell_comb \ramaddr~41 (
// Equation(s):
// \ramaddr~41_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~40_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~40_combout  & ((PC_21))) # (!\ramaddr~40_combout  & (daddr_21))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [21]),
	.datac(\CPU|DP|PCU|PC [21]),
	.datad(\ramaddr~40_combout ),
	.cin(gnd),
	.combout(\ramaddr~41_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~41 .lut_mask = 16'hFA44;
defparam \ramaddr~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N0
cycloneive_lcell_comb \ramaddr~42 (
// Equation(s):
// \ramaddr~42_combout  = (reg_REN1 & (((daddr_20)))) # (!reg_REN1 & ((reg_WEN1 & (daddr_20)) # (!reg_WEN1 & ((PC_20)))))

	.dataa(\CPU|DP|RU|reg_REN~q ),
	.datab(\CPU|DP|RU|reg_WEN~q ),
	.datac(\CPU|CM|daddr [20]),
	.datad(\CPU|DP|PCU|PC [20]),
	.cin(gnd),
	.combout(\ramaddr~42_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~42 .lut_mask = 16'hF1E0;
defparam \ramaddr~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N22
cycloneive_lcell_comb \ramaddr~43 (
// Equation(s):
// \ramaddr~43_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[20]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~42_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[20]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~42_combout ),
	.cin(gnd),
	.combout(\ramaddr~43_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~43 .lut_mask = 16'hDD88;
defparam \ramaddr~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N16
cycloneive_lcell_comb \ramaddr~44 (
// Equation(s):
// \ramaddr~44_combout  = (reg_WEN1 & (((daddr_23)))) # (!reg_WEN1 & ((reg_REN1 & ((daddr_23))) # (!reg_REN1 & (PC_23))))

	.dataa(\CPU|DP|PCU|PC [23]),
	.datab(\CPU|DP|RU|reg_WEN~q ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|CM|daddr [23]),
	.cin(gnd),
	.combout(\ramaddr~44_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~44 .lut_mask = 16'hFE02;
defparam \ramaddr~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N18
cycloneive_lcell_comb \ramaddr~45 (
// Equation(s):
// \ramaddr~45_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[23]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~44_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[23]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~44_combout ),
	.cin(gnd),
	.combout(\ramaddr~45_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~45 .lut_mask = 16'hDD88;
defparam \ramaddr~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N26
cycloneive_lcell_comb \ramaddr~46 (
// Equation(s):
// \ramaddr~46_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[22]~input_o )) # (!\syif.tbCTRL~input_o  & (((reg_REN1) # (reg_WEN1))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[22]~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramaddr~46_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~46 .lut_mask = 16'hDDD8;
defparam \ramaddr~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N12
cycloneive_lcell_comb \ramaddr~47 (
// Equation(s):
// \ramaddr~47_combout  = (\ramaddr~46_combout  & ((\syif.tbCTRL~input_o ) # ((daddr_22)))) # (!\ramaddr~46_combout  & (!\syif.tbCTRL~input_o  & ((PC_22))))

	.dataa(\ramaddr~46_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|CM|daddr [22]),
	.datad(\CPU|DP|PCU|PC [22]),
	.cin(gnd),
	.combout(\ramaddr~47_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~47 .lut_mask = 16'hB9A8;
defparam \ramaddr~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N10
cycloneive_lcell_comb \ramaddr~48 (
// Equation(s):
// \ramaddr~48_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[25]~input_o )) # (!\syif.tbCTRL~input_o  & (((reg_WEN1) # (reg_REN1))))

	.dataa(\syif.addr[25]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RU|reg_WEN~q ),
	.datad(\CPU|DP|RU|reg_REN~q ),
	.cin(gnd),
	.combout(\ramaddr~48_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~48 .lut_mask = 16'hBBB8;
defparam \ramaddr~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N28
cycloneive_lcell_comb \ramaddr~49 (
// Equation(s):
// \ramaddr~49_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~48_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~48_combout  & (daddr_25)) # (!\ramaddr~48_combout  & ((PC_25)))))

	.dataa(\CPU|CM|daddr [25]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|PCU|PC [25]),
	.datad(\ramaddr~48_combout ),
	.cin(gnd),
	.combout(\ramaddr~49_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~49 .lut_mask = 16'hEE30;
defparam \ramaddr~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N0
cycloneive_lcell_comb \ramaddr~50 (
// Equation(s):
// \ramaddr~50_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[24]~input_o )) # (!\syif.tbCTRL~input_o  & (((reg_WEN1) # (reg_REN1))))

	.dataa(\syif.addr[24]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RU|reg_WEN~q ),
	.datad(\CPU|DP|RU|reg_REN~q ),
	.cin(gnd),
	.combout(\ramaddr~50_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~50 .lut_mask = 16'hBBB8;
defparam \ramaddr~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N6
cycloneive_lcell_comb \ramaddr~51 (
// Equation(s):
// \ramaddr~51_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~50_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~50_combout  & (daddr_24)) # (!\ramaddr~50_combout  & ((PC_24)))))

	.dataa(\CPU|CM|daddr [24]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|PCU|PC [24]),
	.datad(\ramaddr~50_combout ),
	.cin(gnd),
	.combout(\ramaddr~51_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~51 .lut_mask = 16'hEE30;
defparam \ramaddr~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N30
cycloneive_lcell_comb \ramaddr~52 (
// Equation(s):
// \ramaddr~52_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[27]~input_o )) # (!\syif.tbCTRL~input_o  & (((!reg_REN1 & !reg_WEN1))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[27]~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramaddr~52_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~52 .lut_mask = 16'h888D;
defparam \ramaddr~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N22
cycloneive_lcell_comb \ramaddr~53 (
// Equation(s):
// \ramaddr~53_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~52_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~52_combout  & (PC_27)) # (!\ramaddr~52_combout  & ((daddr_27)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|PCU|PC [27]),
	.datac(\ramaddr~52_combout ),
	.datad(\CPU|CM|daddr [27]),
	.cin(gnd),
	.combout(\ramaddr~53_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~53 .lut_mask = 16'hE5E0;
defparam \ramaddr~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N10
cycloneive_lcell_comb \ramaddr~54 (
// Equation(s):
// \ramaddr~54_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[26]~input_o )) # (!\syif.tbCTRL~input_o  & (((reg_REN1) # (reg_WEN1))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[26]~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramaddr~54_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~54 .lut_mask = 16'hDDD8;
defparam \ramaddr~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N0
cycloneive_lcell_comb \ramaddr~55 (
// Equation(s):
// \ramaddr~55_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~54_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~54_combout  & ((daddr_26))) # (!\ramaddr~54_combout  & (PC_26))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|PCU|PC [26]),
	.datac(\CPU|CM|daddr [26]),
	.datad(\ramaddr~54_combout ),
	.cin(gnd),
	.combout(\ramaddr~55_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~55 .lut_mask = 16'hFA44;
defparam \ramaddr~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N2
cycloneive_lcell_comb \ramaddr~56 (
// Equation(s):
// \ramaddr~56_combout  = (reg_REN1 & (((daddr_29)))) # (!reg_REN1 & ((reg_WEN1 & ((daddr_29))) # (!reg_WEN1 & (PC_29))))

	.dataa(\CPU|DP|RU|reg_REN~q ),
	.datab(\CPU|DP|RU|reg_WEN~q ),
	.datac(\CPU|DP|PCU|PC [29]),
	.datad(\CPU|CM|daddr [29]),
	.cin(gnd),
	.combout(\ramaddr~56_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~56 .lut_mask = 16'hFE10;
defparam \ramaddr~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N4
cycloneive_lcell_comb \ramaddr~57 (
// Equation(s):
// \ramaddr~57_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[29]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~56_combout )))

	.dataa(\syif.addr[29]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~56_combout ),
	.cin(gnd),
	.combout(\ramaddr~57_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~57 .lut_mask = 16'hBB88;
defparam \ramaddr~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N28
cycloneive_lcell_comb \ramaddr~58 (
// Equation(s):
// \ramaddr~58_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[28]~input_o )) # (!\syif.tbCTRL~input_o  & (((!reg_REN1 & !reg_WEN1))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[28]~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramaddr~58_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~58 .lut_mask = 16'h888D;
defparam \ramaddr~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N10
cycloneive_lcell_comb \ramaddr~59 (
// Equation(s):
// \ramaddr~59_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~58_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~58_combout  & ((PC_28))) # (!\ramaddr~58_combout  & (daddr_28))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [28]),
	.datac(\ramaddr~58_combout ),
	.datad(\CPU|DP|PCU|PC [28]),
	.cin(gnd),
	.combout(\ramaddr~59_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~59 .lut_mask = 16'hF4A4;
defparam \ramaddr~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N12
cycloneive_lcell_comb \ramaddr~60 (
// Equation(s):
// \ramaddr~60_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[31]~input_o )) # (!\syif.tbCTRL~input_o  & (((reg_REN1) # (reg_WEN1))))

	.dataa(\syif.addr[31]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramaddr~60_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~60 .lut_mask = 16'hBBB8;
defparam \ramaddr~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N14
cycloneive_lcell_comb \ramaddr~61 (
// Equation(s):
// \ramaddr~61_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~60_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~60_combout  & (daddr_31)) # (!\ramaddr~60_combout  & ((PC_31)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [31]),
	.datac(\CPU|DP|PCU|PC [31]),
	.datad(\ramaddr~60_combout ),
	.cin(gnd),
	.combout(\ramaddr~61_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~61 .lut_mask = 16'hEE50;
defparam \ramaddr~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N18
cycloneive_lcell_comb \ramaddr~62 (
// Equation(s):
// \ramaddr~62_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[30]~input_o )) # (!\syif.tbCTRL~input_o  & (((!reg_REN1 & !reg_WEN1))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[30]~input_o ),
	.datac(\CPU|DP|RU|reg_REN~q ),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramaddr~62_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~62 .lut_mask = 16'h888D;
defparam \ramaddr~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N0
cycloneive_lcell_comb \ramaddr~63 (
// Equation(s):
// \ramaddr~63_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~62_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~62_combout  & ((PC_30))) # (!\ramaddr~62_combout  & (daddr_30))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [30]),
	.datac(\CPU|DP|PCU|PC [30]),
	.datad(\ramaddr~62_combout ),
	.cin(gnd),
	.combout(\ramaddr~63_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~63 .lut_mask = 16'hFA44;
defparam \ramaddr~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N30
cycloneive_lcell_comb \ramWEN~0 (
// Equation(s):
// \ramWEN~0_combout  = (\syif.tbCTRL~input_o  & (!\syif.WEN~input_o )) # (!\syif.tbCTRL~input_o  & ((!reg_WEN1)))

	.dataa(gnd),
	.datab(\syif.WEN~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramWEN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramWEN~0 .lut_mask = 16'h303F;
defparam \ramWEN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N0
cycloneive_lcell_comb \ramREN~0 (
// Equation(s):
// \ramREN~0_combout  = (\syif.tbCTRL~input_o  & (!\syif.REN~input_o )) # (!\syif.tbCTRL~input_o  & ((reg_WEN1)))

	.dataa(gnd),
	.datab(\syif.REN~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|RU|reg_WEN~q ),
	.cin(gnd),
	.combout(\ramREN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramREN~0 .lut_mask = 16'h3F30;
defparam \ramREN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y72_N19
dffeas CPUCLK(
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\CPUCLK~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\CPUCLK~q ),
	.prn(vcc));
// synopsys translate_off
defparam CPUCLK.is_wysiwyg = "true";
defparam CPUCLK.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N12
cycloneive_lcell_comb \ramstore~0 (
// Equation(s):
// \ramstore~0_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux63))) # (!dcifimemload_20 & (Mux631))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RF|Mux63~23_combout ),
	.datad(\CPU|DP|RF|Mux63~9_combout ),
	.cin(gnd),
	.combout(\ramstore~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~0 .lut_mask = 16'h3210;
defparam \ramstore~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N22
cycloneive_lcell_comb \ramstore~1 (
// Equation(s):
// \ramstore~1_combout  = (\ramstore~0_combout ) # ((\syif.store[0]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[0]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramstore~0_combout ),
	.cin(gnd),
	.combout(\ramstore~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~1 .lut_mask = 16'hFF88;
defparam \ramstore~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N24
cycloneive_lcell_comb \ramstore~2 (
// Equation(s):
// \ramstore~2_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux62)) # (!dcifimemload_20 & ((Mux621)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|RF|Mux62~9_combout ),
	.datad(\CPU|DP|RF|Mux62~21_combout ),
	.cin(gnd),
	.combout(\ramstore~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~2 .lut_mask = 16'h5140;
defparam \ramstore~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N6
cycloneive_lcell_comb \ramstore~3 (
// Equation(s):
// \ramstore~3_combout  = (\ramstore~2_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[1]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[1]~input_o ),
	.datad(\ramstore~2_combout ),
	.cin(gnd),
	.combout(\ramstore~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~3 .lut_mask = 16'hFFA0;
defparam \ramstore~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N2
cycloneive_lcell_comb \ramstore~4 (
// Equation(s):
// \ramstore~4_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux611)) # (!dcifimemload_20 & ((Mux61)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|RF|Mux61~19_combout ),
	.datad(\CPU|DP|RF|Mux61~9_combout ),
	.cin(gnd),
	.combout(\ramstore~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~4 .lut_mask = 16'h5140;
defparam \ramstore~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N20
cycloneive_lcell_comb \ramstore~5 (
// Equation(s):
// \ramstore~5_combout  = (\ramstore~4_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[2]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[2]~input_o ),
	.datac(gnd),
	.datad(\ramstore~4_combout ),
	.cin(gnd),
	.combout(\ramstore~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~5 .lut_mask = 16'hFF88;
defparam \ramstore~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N28
cycloneive_lcell_comb \ramstore~6 (
// Equation(s):
// \ramstore~6_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux60))) # (!dcifimemload_20 & (Mux601))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|RF|Mux60~19_combout ),
	.datad(\CPU|DP|RF|Mux60~9_combout ),
	.cin(gnd),
	.combout(\ramstore~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~6 .lut_mask = 16'h5410;
defparam \ramstore~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N2
cycloneive_lcell_comb \ramstore~7 (
// Equation(s):
// \ramstore~7_combout  = (\ramstore~6_combout ) # ((\syif.store[3]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[3]~input_o ),
	.datab(\ramstore~6_combout ),
	.datac(gnd),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~7 .lut_mask = 16'hEECC;
defparam \ramstore~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N28
cycloneive_lcell_comb \ramstore~8 (
// Equation(s):
// \ramstore~8_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux591)) # (!dcifimemload_20 & ((Mux59)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|RF|Mux59~19_combout ),
	.datad(\CPU|DP|RF|Mux59~9_combout ),
	.cin(gnd),
	.combout(\ramstore~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~8 .lut_mask = 16'h5140;
defparam \ramstore~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N2
cycloneive_lcell_comb \ramstore~9 (
// Equation(s):
// \ramstore~9_combout  = (\ramstore~8_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[4]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[4]~input_o ),
	.datad(\ramstore~8_combout ),
	.cin(gnd),
	.combout(\ramstore~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~9 .lut_mask = 16'hFFA0;
defparam \ramstore~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N20
cycloneive_lcell_comb \ramstore~10 (
// Equation(s):
// \ramstore~10_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux581)) # (!dcifimemload_20 & ((Mux58)))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RF|Mux58~19_combout ),
	.datad(\CPU|DP|RF|Mux58~9_combout ),
	.cin(gnd),
	.combout(\ramstore~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~10 .lut_mask = 16'h3120;
defparam \ramstore~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N22
cycloneive_lcell_comb \ramstore~11 (
// Equation(s):
// \ramstore~11_combout  = (\ramstore~10_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[5]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[5]~input_o ),
	.datad(\ramstore~10_combout ),
	.cin(gnd),
	.combout(\ramstore~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~11 .lut_mask = 16'hFFC0;
defparam \ramstore~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N28
cycloneive_lcell_comb \ramstore~12 (
// Equation(s):
// \ramstore~12_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux571)) # (!dcifimemload_20 & ((Mux57)))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RF|Mux57~19_combout ),
	.datad(\CPU|DP|RF|Mux57~9_combout ),
	.cin(gnd),
	.combout(\ramstore~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~12 .lut_mask = 16'h3120;
defparam \ramstore~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N6
cycloneive_lcell_comb \ramstore~13 (
// Equation(s):
// \ramstore~13_combout  = (\ramstore~12_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[6]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[6]~input_o ),
	.datad(\ramstore~12_combout ),
	.cin(gnd),
	.combout(\ramstore~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~13 .lut_mask = 16'hFFC0;
defparam \ramstore~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N12
cycloneive_lcell_comb \ramstore~14 (
// Equation(s):
// \ramstore~14_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux561)) # (!dcifimemload_20 & ((Mux56)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|RF|Mux56~19_combout ),
	.datad(\CPU|DP|RF|Mux56~9_combout ),
	.cin(gnd),
	.combout(\ramstore~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~14 .lut_mask = 16'h5140;
defparam \ramstore~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N6
cycloneive_lcell_comb \ramstore~15 (
// Equation(s):
// \ramstore~15_combout  = (\ramstore~14_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[7]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[7]~input_o ),
	.datac(gnd),
	.datad(\ramstore~14_combout ),
	.cin(gnd),
	.combout(\ramstore~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~15 .lut_mask = 16'hFF88;
defparam \ramstore~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N28
cycloneive_lcell_comb \ramstore~16 (
// Equation(s):
// \ramstore~16_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux551))) # (!dcifimemload_20 & (Mux55))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|RF|Mux55~9_combout ),
	.datac(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datad(\CPU|DP|RF|Mux55~19_combout ),
	.cin(gnd),
	.combout(\ramstore~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~16 .lut_mask = 16'h5404;
defparam \ramstore~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N18
cycloneive_lcell_comb \ramstore~17 (
// Equation(s):
// \ramstore~17_combout  = (\ramstore~16_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[8]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[8]~input_o ),
	.datac(gnd),
	.datad(\ramstore~16_combout ),
	.cin(gnd),
	.combout(\ramstore~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~17 .lut_mask = 16'hFF88;
defparam \ramstore~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N0
cycloneive_lcell_comb \ramstore~18 (
// Equation(s):
// \ramstore~18_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux541))) # (!dcifimemload_20 & (Mux54))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|RF|Mux54~9_combout ),
	.datac(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datad(\CPU|DP|RF|Mux54~19_combout ),
	.cin(gnd),
	.combout(\ramstore~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~18 .lut_mask = 16'h5404;
defparam \ramstore~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N6
cycloneive_lcell_comb \ramstore~19 (
// Equation(s):
// \ramstore~19_combout  = (\ramstore~18_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[9]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[9]~input_o ),
	.datad(\ramstore~18_combout ),
	.cin(gnd),
	.combout(\ramstore~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~19 .lut_mask = 16'hFFA0;
defparam \ramstore~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N24
cycloneive_lcell_comb \ramstore~20 (
// Equation(s):
// \ramstore~20_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux531))) # (!dcifimemload_20 & (Mux53))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|RF|Mux53~9_combout ),
	.datac(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datad(\CPU|DP|RF|Mux53~19_combout ),
	.cin(gnd),
	.combout(\ramstore~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~20 .lut_mask = 16'h5404;
defparam \ramstore~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N22
cycloneive_lcell_comb \ramstore~21 (
// Equation(s):
// \ramstore~21_combout  = (\ramstore~20_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[10]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[10]~input_o ),
	.datad(\ramstore~20_combout ),
	.cin(gnd),
	.combout(\ramstore~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~21 .lut_mask = 16'hFFC0;
defparam \ramstore~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N12
cycloneive_lcell_comb \ramstore~22 (
// Equation(s):
// \ramstore~22_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux521))) # (!dcifimemload_20 & (Mux52))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|RF|Mux52~9_combout ),
	.datac(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datad(\CPU|DP|RF|Mux52~19_combout ),
	.cin(gnd),
	.combout(\ramstore~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~22 .lut_mask = 16'h5404;
defparam \ramstore~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N2
cycloneive_lcell_comb \ramstore~23 (
// Equation(s):
// \ramstore~23_combout  = (\ramstore~22_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[11]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[11]~input_o ),
	.datad(\ramstore~22_combout ),
	.cin(gnd),
	.combout(\ramstore~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~23 .lut_mask = 16'hFFC0;
defparam \ramstore~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N28
cycloneive_lcell_comb \ramstore~24 (
// Equation(s):
// \ramstore~24_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux511))) # (!dcifimemload_20 & (Mux51))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|RF|Mux51~9_combout ),
	.datac(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datad(\CPU|DP|RF|Mux51~19_combout ),
	.cin(gnd),
	.combout(\ramstore~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~24 .lut_mask = 16'h5404;
defparam \ramstore~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N22
cycloneive_lcell_comb \ramstore~25 (
// Equation(s):
// \ramstore~25_combout  = (\ramstore~24_combout ) # ((\syif.store[12]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[12]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramstore~24_combout ),
	.cin(gnd),
	.combout(\ramstore~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~25 .lut_mask = 16'hFF88;
defparam \ramstore~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N12
cycloneive_lcell_comb \ramstore~26 (
// Equation(s):
// \ramstore~26_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux501)) # (!dcifimemload_20 & ((Mux50)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|RF|Mux50~19_combout ),
	.datad(\CPU|DP|RF|Mux50~9_combout ),
	.cin(gnd),
	.combout(\ramstore~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~26 .lut_mask = 16'h5140;
defparam \ramstore~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N6
cycloneive_lcell_comb \ramstore~27 (
// Equation(s):
// \ramstore~27_combout  = (\ramstore~26_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[13]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[13]~input_o ),
	.datad(\ramstore~26_combout ),
	.cin(gnd),
	.combout(\ramstore~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~27 .lut_mask = 16'hFFC0;
defparam \ramstore~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N12
cycloneive_lcell_comb \ramstore~28 (
// Equation(s):
// \ramstore~28_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux491)) # (!dcifimemload_20 & ((Mux49)))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RF|Mux49~19_combout ),
	.datad(\CPU|DP|RF|Mux49~9_combout ),
	.cin(gnd),
	.combout(\ramstore~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~28 .lut_mask = 16'h3120;
defparam \ramstore~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N18
cycloneive_lcell_comb \ramstore~29 (
// Equation(s):
// \ramstore~29_combout  = (\ramstore~28_combout ) # ((\syif.store[14]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[14]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramstore~28_combout ),
	.cin(gnd),
	.combout(\ramstore~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~29 .lut_mask = 16'hFF88;
defparam \ramstore~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N0
cycloneive_lcell_comb \ramstore~30 (
// Equation(s):
// \ramstore~30_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux481)) # (!dcifimemload_20 & ((Mux48)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|RF|Mux48~19_combout ),
	.datad(\CPU|DP|RF|Mux48~9_combout ),
	.cin(gnd),
	.combout(\ramstore~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~30 .lut_mask = 16'h5140;
defparam \ramstore~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N26
cycloneive_lcell_comb \ramstore~31 (
// Equation(s):
// \ramstore~31_combout  = (\ramstore~30_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[15]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[15]~input_o ),
	.datad(\ramstore~30_combout ),
	.cin(gnd),
	.combout(\ramstore~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~31 .lut_mask = 16'hFFA0;
defparam \ramstore~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N24
cycloneive_lcell_comb \ramstore~32 (
// Equation(s):
// \ramstore~32_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux471)) # (!dcifimemload_20 & ((Mux47)))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RF|Mux47~19_combout ),
	.datad(\CPU|DP|RF|Mux47~9_combout ),
	.cin(gnd),
	.combout(\ramstore~32_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~32 .lut_mask = 16'h3120;
defparam \ramstore~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N22
cycloneive_lcell_comb \ramstore~33 (
// Equation(s):
// \ramstore~33_combout  = (\ramstore~32_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[16]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[16]~input_o ),
	.datad(\ramstore~32_combout ),
	.cin(gnd),
	.combout(\ramstore~33_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~33 .lut_mask = 16'hFFC0;
defparam \ramstore~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N20
cycloneive_lcell_comb \ramstore~34 (
// Equation(s):
// \ramstore~34_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux461))) # (!dcifimemload_20 & (Mux46))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|RF|Mux46~9_combout ),
	.datac(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datad(\CPU|DP|RF|Mux46~19_combout ),
	.cin(gnd),
	.combout(\ramstore~34_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~34 .lut_mask = 16'h5404;
defparam \ramstore~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N2
cycloneive_lcell_comb \ramstore~35 (
// Equation(s):
// \ramstore~35_combout  = (\ramstore~34_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[17]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[17]~input_o ),
	.datac(gnd),
	.datad(\ramstore~34_combout ),
	.cin(gnd),
	.combout(\ramstore~35_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~35 .lut_mask = 16'hFF88;
defparam \ramstore~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N20
cycloneive_lcell_comb \ramstore~36 (
// Equation(s):
// \ramstore~36_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux451))) # (!dcifimemload_20 & (Mux45))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|RF|Mux45~9_combout ),
	.datad(\CPU|DP|RF|Mux45~19_combout ),
	.cin(gnd),
	.combout(\ramstore~36_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~36 .lut_mask = 16'h5410;
defparam \ramstore~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N14
cycloneive_lcell_comb \ramstore~37 (
// Equation(s):
// \ramstore~37_combout  = (\ramstore~36_combout ) # ((\syif.store[18]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[18]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~36_combout ),
	.cin(gnd),
	.combout(\ramstore~37_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~37 .lut_mask = 16'hFFA0;
defparam \ramstore~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N0
cycloneive_lcell_comb \ramstore~38 (
// Equation(s):
// \ramstore~38_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux441)) # (!dcifimemload_20 & ((Mux44)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|RF|Mux44~19_combout ),
	.datac(\CPU|DP|RF|Mux44~9_combout ),
	.datad(\CPU|CM|dcif.imemload[20]~10_combout ),
	.cin(gnd),
	.combout(\ramstore~38_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~38 .lut_mask = 16'h4450;
defparam \ramstore~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N22
cycloneive_lcell_comb \ramstore~39 (
// Equation(s):
// \ramstore~39_combout  = (\ramstore~38_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[19]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[19]~input_o ),
	.datad(\ramstore~38_combout ),
	.cin(gnd),
	.combout(\ramstore~39_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~39 .lut_mask = 16'hFFA0;
defparam \ramstore~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N24
cycloneive_lcell_comb \ramstore~40 (
// Equation(s):
// \ramstore~40_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux431))) # (!dcifimemload_20 & (Mux43))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|RF|Mux43~9_combout ),
	.datad(\CPU|DP|RF|Mux43~19_combout ),
	.cin(gnd),
	.combout(\ramstore~40_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~40 .lut_mask = 16'h5410;
defparam \ramstore~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N14
cycloneive_lcell_comb \ramstore~41 (
// Equation(s):
// \ramstore~41_combout  = (\ramstore~40_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[20]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\ramstore~40_combout ),
	.datac(gnd),
	.datad(\syif.store[20]~input_o ),
	.cin(gnd),
	.combout(\ramstore~41_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~41 .lut_mask = 16'hEECC;
defparam \ramstore~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N10
cycloneive_lcell_comb \ramstore~42 (
// Equation(s):
// \ramstore~42_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux421)) # (!dcifimemload_20 & ((Mux42)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|RF|Mux42~19_combout ),
	.datad(\CPU|DP|RF|Mux42~9_combout ),
	.cin(gnd),
	.combout(\ramstore~42_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~42 .lut_mask = 16'h5140;
defparam \ramstore~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N4
cycloneive_lcell_comb \ramstore~43 (
// Equation(s):
// \ramstore~43_combout  = (\ramstore~42_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[21]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[21]~input_o ),
	.datac(gnd),
	.datad(\ramstore~42_combout ),
	.cin(gnd),
	.combout(\ramstore~43_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~43 .lut_mask = 16'hFF88;
defparam \ramstore~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N0
cycloneive_lcell_comb \ramstore~44 (
// Equation(s):
// \ramstore~44_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux411))) # (!dcifimemload_20 & (Mux41))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|RF|Mux41~9_combout ),
	.datad(\CPU|DP|RF|Mux41~19_combout ),
	.cin(gnd),
	.combout(\ramstore~44_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~44 .lut_mask = 16'h5410;
defparam \ramstore~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N2
cycloneive_lcell_comb \ramstore~45 (
// Equation(s):
// \ramstore~45_combout  = (\ramstore~44_combout ) # ((\syif.store[22]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[22]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~44_combout ),
	.cin(gnd),
	.combout(\ramstore~45_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~45 .lut_mask = 16'hFFC0;
defparam \ramstore~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N0
cycloneive_lcell_comb \ramstore~46 (
// Equation(s):
// \ramstore~46_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux401))) # (!dcifimemload_20 & (Mux40))))

	.dataa(\CPU|DP|RF|Mux40~9_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RF|Mux40~19_combout ),
	.datad(\CPU|CM|dcif.imemload[20]~10_combout ),
	.cin(gnd),
	.combout(\ramstore~46_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~46 .lut_mask = 16'h3022;
defparam \ramstore~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N2
cycloneive_lcell_comb \ramstore~47 (
// Equation(s):
// \ramstore~47_combout  = (\ramstore~46_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[23]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[23]~input_o ),
	.datad(\ramstore~46_combout ),
	.cin(gnd),
	.combout(\ramstore~47_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~47 .lut_mask = 16'hFFC0;
defparam \ramstore~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N24
cycloneive_lcell_comb \ramstore~48 (
// Equation(s):
// \ramstore~48_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux391))) # (!dcifimemload_20 & (Mux39))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RF|Mux39~9_combout ),
	.datad(\CPU|DP|RF|Mux39~19_combout ),
	.cin(gnd),
	.combout(\ramstore~48_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~48 .lut_mask = 16'h3210;
defparam \ramstore~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N14
cycloneive_lcell_comb \ramstore~49 (
// Equation(s):
// \ramstore~49_combout  = (\ramstore~48_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[24]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[24]~input_o ),
	.datac(gnd),
	.datad(\ramstore~48_combout ),
	.cin(gnd),
	.combout(\ramstore~49_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~49 .lut_mask = 16'hFF88;
defparam \ramstore~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N14
cycloneive_lcell_comb \ramstore~50 (
// Equation(s):
// \ramstore~50_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux381)) # (!dcifimemload_20 & ((Mux38)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|RF|Mux38~19_combout ),
	.datad(\CPU|DP|RF|Mux38~9_combout ),
	.cin(gnd),
	.combout(\ramstore~50_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~50 .lut_mask = 16'h5140;
defparam \ramstore~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N28
cycloneive_lcell_comb \ramstore~51 (
// Equation(s):
// \ramstore~51_combout  = (\ramstore~50_combout ) # ((\syif.store[25]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[25]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~50_combout ),
	.cin(gnd),
	.combout(\ramstore~51_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~51 .lut_mask = 16'hFFC0;
defparam \ramstore~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N28
cycloneive_lcell_comb \ramstore~52 (
// Equation(s):
// \ramstore~52_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux371))) # (!dcifimemload_20 & (Mux37))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|RF|Mux37~9_combout ),
	.datac(\CPU|DP|RF|Mux37~19_combout ),
	.datad(\CPU|CM|dcif.imemload[20]~10_combout ),
	.cin(gnd),
	.combout(\ramstore~52_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~52 .lut_mask = 16'h5044;
defparam \ramstore~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N18
cycloneive_lcell_comb \ramstore~53 (
// Equation(s):
// \ramstore~53_combout  = (\ramstore~52_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[26]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[26]~input_o ),
	.datac(gnd),
	.datad(\ramstore~52_combout ),
	.cin(gnd),
	.combout(\ramstore~53_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~53 .lut_mask = 16'hFF88;
defparam \ramstore~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N4
cycloneive_lcell_comb \ramstore~54 (
// Equation(s):
// \ramstore~54_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux361)) # (!dcifimemload_20 & ((Mux36)))))

	.dataa(\CPU|DP|RF|Mux36~19_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datad(\CPU|DP|RF|Mux36~9_combout ),
	.cin(gnd),
	.combout(\ramstore~54_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~54 .lut_mask = 16'h2320;
defparam \ramstore~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N2
cycloneive_lcell_comb \ramstore~55 (
// Equation(s):
// \ramstore~55_combout  = (\ramstore~54_combout ) # ((\syif.store[27]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[27]~input_o ),
	.datac(\ramstore~54_combout ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~55_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~55 .lut_mask = 16'hFCF0;
defparam \ramstore~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N16
cycloneive_lcell_comb \ramstore~56 (
// Equation(s):
// \ramstore~56_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux351)) # (!dcifimemload_20 & ((Mux35)))))

	.dataa(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|RF|Mux35~19_combout ),
	.datad(\CPU|DP|RF|Mux35~9_combout ),
	.cin(gnd),
	.combout(\ramstore~56_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~56 .lut_mask = 16'h3120;
defparam \ramstore~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N10
cycloneive_lcell_comb \ramstore~57 (
// Equation(s):
// \ramstore~57_combout  = (\ramstore~56_combout ) # ((\syif.store[28]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[28]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramstore~56_combout ),
	.cin(gnd),
	.combout(\ramstore~57_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~57 .lut_mask = 16'hFF88;
defparam \ramstore~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N0
cycloneive_lcell_comb \ramstore~58 (
// Equation(s):
// \ramstore~58_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux341)) # (!dcifimemload_20 & ((Mux34)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|RF|Mux34~19_combout ),
	.datad(\CPU|DP|RF|Mux34~9_combout ),
	.cin(gnd),
	.combout(\ramstore~58_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~58 .lut_mask = 16'h5140;
defparam \ramstore~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N2
cycloneive_lcell_comb \ramstore~59 (
// Equation(s):
// \ramstore~59_combout  = (\ramstore~58_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[29]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[29]~input_o ),
	.datad(\ramstore~58_combout ),
	.cin(gnd),
	.combout(\ramstore~59_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~59 .lut_mask = 16'hFFA0;
defparam \ramstore~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N12
cycloneive_lcell_comb \ramstore~60 (
// Equation(s):
// \ramstore~60_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & ((Mux331))) # (!dcifimemload_20 & (Mux33))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datac(\CPU|DP|RF|Mux33~9_combout ),
	.datad(\CPU|DP|RF|Mux33~19_combout ),
	.cin(gnd),
	.combout(\ramstore~60_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~60 .lut_mask = 16'h5410;
defparam \ramstore~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N26
cycloneive_lcell_comb \ramstore~61 (
// Equation(s):
// \ramstore~61_combout  = (\ramstore~60_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[30]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[30]~input_o ),
	.datad(\ramstore~60_combout ),
	.cin(gnd),
	.combout(\ramstore~61_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~61 .lut_mask = 16'hFFA0;
defparam \ramstore~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N8
cycloneive_lcell_comb \ramstore~62 (
// Equation(s):
// \ramstore~62_combout  = (!\syif.tbCTRL~input_o  & ((dcifimemload_20 & (Mux321)) # (!dcifimemload_20 & ((Mux32)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|RF|Mux32~19_combout ),
	.datac(\CPU|CM|dcif.imemload[20]~10_combout ),
	.datad(\CPU|DP|RF|Mux32~9_combout ),
	.cin(gnd),
	.combout(\ramstore~62_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~62 .lut_mask = 16'h4540;
defparam \ramstore~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N6
cycloneive_lcell_comb \ramstore~63 (
// Equation(s):
// \ramstore~63_combout  = (\ramstore~62_combout ) # ((\syif.store[31]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[31]~input_o ),
	.datab(gnd),
	.datac(\ramstore~62_combout ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~63_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~63 .lut_mask = 16'hFAF0;
defparam \ramstore~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y72_N1
dffeas \count[3] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[3]~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[3]),
	.prn(vcc));
// synopsys translate_off
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y72_N5
dffeas \count[2] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[2]~1_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[2]),
	.prn(vcc));
// synopsys translate_off
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y72_N13
dffeas \count[1] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[1]~2_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[1]),
	.prn(vcc));
// synopsys translate_off
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y72_N9
dffeas \count[0] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[0]),
	.prn(vcc));
// synopsys translate_off
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y72_N10
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (!count[1] & (!count[2] & (!count[0] & !count[3])))

	.dataa(count[1]),
	.datab(count[2]),
	.datac(count[0]),
	.datad(count[3]),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h0001;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y72_N18
cycloneive_lcell_comb \CPUCLK~0 (
// Equation(s):
// \CPUCLK~0_combout  = \CPUCLK~q  $ (\Equal0~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\CPUCLK~q ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\CPUCLK~0_combout ),
	.cout());
// synopsys translate_off
defparam \CPUCLK~0 .lut_mask = 16'h0FF0;
defparam \CPUCLK~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y72_N0
cycloneive_lcell_comb \count[3]~0 (
// Equation(s):
// \count[3]~0_combout  = count[3] $ (((count[1] & (count[0] & count[2]))))

	.dataa(count[1]),
	.datab(count[0]),
	.datac(count[3]),
	.datad(count[2]),
	.cin(gnd),
	.combout(\count[3]~0_combout ),
	.cout());
// synopsys translate_off
defparam \count[3]~0 .lut_mask = 16'h78F0;
defparam \count[3]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y72_N4
cycloneive_lcell_comb \count[2]~1 (
// Equation(s):
// \count[2]~1_combout  = count[2] $ (((count[0] & count[1])))

	.dataa(gnd),
	.datab(count[0]),
	.datac(count[2]),
	.datad(count[1]),
	.cin(gnd),
	.combout(\count[2]~1_combout ),
	.cout());
// synopsys translate_off
defparam \count[2]~1 .lut_mask = 16'h3CF0;
defparam \count[2]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y72_N12
cycloneive_lcell_comb \count[1]~2 (
// Equation(s):
// \count[1]~2_combout  = count[0] $ (count[1])

	.dataa(gnd),
	.datab(count[0]),
	.datac(count[1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \count[1]~2 .lut_mask = 16'h3C3C;
defparam \count[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y72_N8
cycloneive_lcell_comb \count~3 (
// Equation(s):
// \count~3_combout  = (!count[0] & ((count[1]) # ((count[2]) # (count[3]))))

	.dataa(count[1]),
	.datab(count[2]),
	.datac(count[0]),
	.datad(count[3]),
	.cin(gnd),
	.combout(\count~3_combout ),
	.cout());
// synopsys translate_off
defparam \count~3 .lut_mask = 16'h0F0E;
defparam \count~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N26
cycloneive_lcell_comb \ramaddr~29_wirecell (
// Equation(s):
// \ramaddr~29_wirecell_combout  = !\ramaddr~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\ramaddr~29_combout ),
	.cin(gnd),
	.combout(\ramaddr~29_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29_wirecell .lut_mask = 16'h00FF;
defparam \ramaddr~29_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: JTAG_X1_Y37_N0
cycloneive_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

// Location: FF_X36_Y39_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~10 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11 .lut_mask = 16'h5AAF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X43_Y41_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y41_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y41_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y41_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y41_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X39_Y41_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y40_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .lut_mask = 16'hFA50;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y40_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .lut_mask = 16'hAAB0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y40_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .lut_mask = 16'hFAAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y41_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .lut_mask = 16'hF780;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .lut_mask = 16'h020A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .lut_mask = 16'hAAE0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .lut_mask = 16'hBA10;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y40_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .lut_mask = 16'h0004;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y39_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .lut_mask = 16'h0400;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y39_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 .lut_mask = 16'h5488;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .lut_mask = 16'h4F41;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .lut_mask = 16'h5000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y40_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .lut_mask = 16'h1AF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .lut_mask = 16'hFF01;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .lut_mask = 16'h0004;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y40_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .lut_mask = 16'hF0F8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .lut_mask = 16'h0504;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .lut_mask = 16'h00EC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 .lut_mask = 16'h0CAE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .lut_mask = 16'h2D8B;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .lut_mask = 16'h5090;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N8
cycloneive_io_ibuf \syif.tbCTRL~input (
	.i(\syif.tbCTRL ),
	.ibar(gnd),
	.o(\syif.tbCTRL~input_o ));
// synopsys translate_off
defparam \syif.tbCTRL~input .bus_hold = "false";
defparam \syif.tbCTRL~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N1
cycloneive_io_ibuf \syif.addr[1]~input (
	.i(\syif.addr [1]),
	.ibar(gnd),
	.o(\syif.addr[1]~input_o ));
// synopsys translate_off
defparam \syif.addr[1]~input .bus_hold = "false";
defparam \syif.addr[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y0_N1
cycloneive_io_ibuf \syif.addr[0]~input (
	.i(\syif.addr [0]),
	.ibar(gnd),
	.o(\syif.addr[0]~input_o ));
// synopsys translate_off
defparam \syif.addr[0]~input .bus_hold = "false";
defparam \syif.addr[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N8
cycloneive_io_ibuf \syif.addr[3]~input (
	.i(\syif.addr [3]),
	.ibar(gnd),
	.o(\syif.addr[3]~input_o ));
// synopsys translate_off
defparam \syif.addr[3]~input .bus_hold = "false";
defparam \syif.addr[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y31_N8
cycloneive_io_ibuf \syif.addr[2]~input (
	.i(\syif.addr [2]),
	.ibar(gnd),
	.o(\syif.addr[2]~input_o ));
// synopsys translate_off
defparam \syif.addr[2]~input .bus_hold = "false";
defparam \syif.addr[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N8
cycloneive_io_ibuf \syif.addr[5]~input (
	.i(\syif.addr [5]),
	.ibar(gnd),
	.o(\syif.addr[5]~input_o ));
// synopsys translate_off
defparam \syif.addr[5]~input .bus_hold = "false";
defparam \syif.addr[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y73_N15
cycloneive_io_ibuf \syif.addr[4]~input (
	.i(\syif.addr [4]),
	.ibar(gnd),
	.o(\syif.addr[4]~input_o ));
// synopsys translate_off
defparam \syif.addr[4]~input .bus_hold = "false";
defparam \syif.addr[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N1
cycloneive_io_ibuf \syif.addr[7]~input (
	.i(\syif.addr [7]),
	.ibar(gnd),
	.o(\syif.addr[7]~input_o ));
// synopsys translate_off
defparam \syif.addr[7]~input .bus_hold = "false";
defparam \syif.addr[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N22
cycloneive_io_ibuf \syif.addr[6]~input (
	.i(\syif.addr [6]),
	.ibar(gnd),
	.o(\syif.addr[6]~input_o ));
// synopsys translate_off
defparam \syif.addr[6]~input .bus_hold = "false";
defparam \syif.addr[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N22
cycloneive_io_ibuf \syif.addr[9]~input (
	.i(\syif.addr [9]),
	.ibar(gnd),
	.o(\syif.addr[9]~input_o ));
// synopsys translate_off
defparam \syif.addr[9]~input .bus_hold = "false";
defparam \syif.addr[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N8
cycloneive_io_ibuf \syif.addr[8]~input (
	.i(\syif.addr [8]),
	.ibar(gnd),
	.o(\syif.addr[8]~input_o ));
// synopsys translate_off
defparam \syif.addr[8]~input .bus_hold = "false";
defparam \syif.addr[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y32_N15
cycloneive_io_ibuf \syif.addr[11]~input (
	.i(\syif.addr [11]),
	.ibar(gnd),
	.o(\syif.addr[11]~input_o ));
// synopsys translate_off
defparam \syif.addr[11]~input .bus_hold = "false";
defparam \syif.addr[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N15
cycloneive_io_ibuf \syif.addr[10]~input (
	.i(\syif.addr [10]),
	.ibar(gnd),
	.o(\syif.addr[10]~input_o ));
// synopsys translate_off
defparam \syif.addr[10]~input .bus_hold = "false";
defparam \syif.addr[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y35_N15
cycloneive_io_ibuf \syif.addr[13]~input (
	.i(\syif.addr [13]),
	.ibar(gnd),
	.o(\syif.addr[13]~input_o ));
// synopsys translate_off
defparam \syif.addr[13]~input .bus_hold = "false";
defparam \syif.addr[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N22
cycloneive_io_ibuf \syif.addr[12]~input (
	.i(\syif.addr [12]),
	.ibar(gnd),
	.o(\syif.addr[12]~input_o ));
// synopsys translate_off
defparam \syif.addr[12]~input .bus_hold = "false";
defparam \syif.addr[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N8
cycloneive_io_ibuf \syif.addr[15]~input (
	.i(\syif.addr [15]),
	.ibar(gnd),
	.o(\syif.addr[15]~input_o ));
// synopsys translate_off
defparam \syif.addr[15]~input .bus_hold = "false";
defparam \syif.addr[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N22
cycloneive_io_ibuf \syif.addr[14]~input (
	.i(\syif.addr [14]),
	.ibar(gnd),
	.o(\syif.addr[14]~input_o ));
// synopsys translate_off
defparam \syif.addr[14]~input .bus_hold = "false";
defparam \syif.addr[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y73_N22
cycloneive_io_ibuf \syif.addr[17]~input (
	.i(\syif.addr [17]),
	.ibar(gnd),
	.o(\syif.addr[17]~input_o ));
// synopsys translate_off
defparam \syif.addr[17]~input .bus_hold = "false";
defparam \syif.addr[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y73_N1
cycloneive_io_ibuf \syif.addr[16]~input (
	.i(\syif.addr [16]),
	.ibar(gnd),
	.o(\syif.addr[16]~input_o ));
// synopsys translate_off
defparam \syif.addr[16]~input .bus_hold = "false";
defparam \syif.addr[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N8
cycloneive_io_ibuf \syif.addr[19]~input (
	.i(\syif.addr [19]),
	.ibar(gnd),
	.o(\syif.addr[19]~input_o ));
// synopsys translate_off
defparam \syif.addr[19]~input .bus_hold = "false";
defparam \syif.addr[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N22
cycloneive_io_ibuf \syif.addr[18]~input (
	.i(\syif.addr [18]),
	.ibar(gnd),
	.o(\syif.addr[18]~input_o ));
// synopsys translate_off
defparam \syif.addr[18]~input .bus_hold = "false";
defparam \syif.addr[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N1
cycloneive_io_ibuf \syif.addr[21]~input (
	.i(\syif.addr [21]),
	.ibar(gnd),
	.o(\syif.addr[21]~input_o ));
// synopsys translate_off
defparam \syif.addr[21]~input .bus_hold = "false";
defparam \syif.addr[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N15
cycloneive_io_ibuf \syif.addr[20]~input (
	.i(\syif.addr [20]),
	.ibar(gnd),
	.o(\syif.addr[20]~input_o ));
// synopsys translate_off
defparam \syif.addr[20]~input .bus_hold = "false";
defparam \syif.addr[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N8
cycloneive_io_ibuf \syif.addr[23]~input (
	.i(\syif.addr [23]),
	.ibar(gnd),
	.o(\syif.addr[23]~input_o ));
// synopsys translate_off
defparam \syif.addr[23]~input .bus_hold = "false";
defparam \syif.addr[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N8
cycloneive_io_ibuf \syif.addr[22]~input (
	.i(\syif.addr [22]),
	.ibar(gnd),
	.o(\syif.addr[22]~input_o ));
// synopsys translate_off
defparam \syif.addr[22]~input .bus_hold = "false";
defparam \syif.addr[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N15
cycloneive_io_ibuf \syif.addr[25]~input (
	.i(\syif.addr [25]),
	.ibar(gnd),
	.o(\syif.addr[25]~input_o ));
// synopsys translate_off
defparam \syif.addr[25]~input .bus_hold = "false";
defparam \syif.addr[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N8
cycloneive_io_ibuf \syif.addr[24]~input (
	.i(\syif.addr [24]),
	.ibar(gnd),
	.o(\syif.addr[24]~input_o ));
// synopsys translate_off
defparam \syif.addr[24]~input .bus_hold = "false";
defparam \syif.addr[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X79_Y73_N1
cycloneive_io_ibuf \syif.addr[27]~input (
	.i(\syif.addr [27]),
	.ibar(gnd),
	.o(\syif.addr[27]~input_o ));
// synopsys translate_off
defparam \syif.addr[27]~input .bus_hold = "false";
defparam \syif.addr[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N15
cycloneive_io_ibuf \syif.addr[26]~input (
	.i(\syif.addr [26]),
	.ibar(gnd),
	.o(\syif.addr[26]~input_o ));
// synopsys translate_off
defparam \syif.addr[26]~input .bus_hold = "false";
defparam \syif.addr[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N22
cycloneive_io_ibuf \syif.addr[29]~input (
	.i(\syif.addr [29]),
	.ibar(gnd),
	.o(\syif.addr[29]~input_o ));
// synopsys translate_off
defparam \syif.addr[29]~input .bus_hold = "false";
defparam \syif.addr[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N1
cycloneive_io_ibuf \syif.addr[28]~input (
	.i(\syif.addr [28]),
	.ibar(gnd),
	.o(\syif.addr[28]~input_o ));
// synopsys translate_off
defparam \syif.addr[28]~input .bus_hold = "false";
defparam \syif.addr[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N22
cycloneive_io_ibuf \syif.addr[31]~input (
	.i(\syif.addr [31]),
	.ibar(gnd),
	.o(\syif.addr[31]~input_o ));
// synopsys translate_off
defparam \syif.addr[31]~input .bus_hold = "false";
defparam \syif.addr[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y33_N8
cycloneive_io_ibuf \syif.addr[30]~input (
	.i(\syif.addr [30]),
	.ibar(gnd),
	.o(\syif.addr[30]~input_o ));
// synopsys translate_off
defparam \syif.addr[30]~input .bus_hold = "false";
defparam \syif.addr[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y34_N15
cycloneive_io_ibuf \syif.WEN~input (
	.i(\syif.WEN ),
	.ibar(gnd),
	.o(\syif.WEN~input_o ));
// synopsys translate_off
defparam \syif.WEN~input .bus_hold = "false";
defparam \syif.WEN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N1
cycloneive_io_ibuf \syif.REN~input (
	.i(\syif.REN ),
	.ibar(gnd),
	.o(\syif.REN~input_o ));
// synopsys translate_off
defparam \syif.REN~input .bus_hold = "false";
defparam \syif.REN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N15
cycloneive_io_ibuf \nRST~input (
	.i(nRST),
	.ibar(gnd),
	.o(\nRST~input_o ));
// synopsys translate_off
defparam \nRST~input .bus_hold = "false";
defparam \nRST~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N8
cycloneive_io_ibuf \CLK~input (
	.i(CLK),
	.ibar(gnd),
	.o(\CLK~input_o ));
// synopsys translate_off
defparam \CLK~input .bus_hold = "false";
defparam \CLK~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y73_N22
cycloneive_io_ibuf \syif.store[0]~input (
	.i(\syif.store [0]),
	.ibar(gnd),
	.o(\syif.store[0]~input_o ));
// synopsys translate_off
defparam \syif.store[0]~input .bus_hold = "false";
defparam \syif.store[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N1
cycloneive_io_ibuf \syif.store[1]~input (
	.i(\syif.store [1]),
	.ibar(gnd),
	.o(\syif.store[1]~input_o ));
// synopsys translate_off
defparam \syif.store[1]~input .bus_hold = "false";
defparam \syif.store[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y73_N15
cycloneive_io_ibuf \syif.store[2]~input (
	.i(\syif.store [2]),
	.ibar(gnd),
	.o(\syif.store[2]~input_o ));
// synopsys translate_off
defparam \syif.store[2]~input .bus_hold = "false";
defparam \syif.store[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y35_N22
cycloneive_io_ibuf \syif.store[3]~input (
	.i(\syif.store [3]),
	.ibar(gnd),
	.o(\syif.store[3]~input_o ));
// synopsys translate_off
defparam \syif.store[3]~input .bus_hold = "false";
defparam \syif.store[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N15
cycloneive_io_ibuf \syif.store[4]~input (
	.i(\syif.store [4]),
	.ibar(gnd),
	.o(\syif.store[4]~input_o ));
// synopsys translate_off
defparam \syif.store[4]~input .bus_hold = "false";
defparam \syif.store[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y0_N15
cycloneive_io_ibuf \syif.store[5]~input (
	.i(\syif.store [5]),
	.ibar(gnd),
	.o(\syif.store[5]~input_o ));
// synopsys translate_off
defparam \syif.store[5]~input .bus_hold = "false";
defparam \syif.store[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N8
cycloneive_io_ibuf \syif.store[6]~input (
	.i(\syif.store [6]),
	.ibar(gnd),
	.o(\syif.store[6]~input_o ));
// synopsys translate_off
defparam \syif.store[6]~input .bus_hold = "false";
defparam \syif.store[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N8
cycloneive_io_ibuf \syif.store[7]~input (
	.i(\syif.store [7]),
	.ibar(gnd),
	.o(\syif.store[7]~input_o ));
// synopsys translate_off
defparam \syif.store[7]~input .bus_hold = "false";
defparam \syif.store[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y73_N1
cycloneive_io_ibuf \syif.store[8]~input (
	.i(\syif.store [8]),
	.ibar(gnd),
	.o(\syif.store[8]~input_o ));
// synopsys translate_off
defparam \syif.store[8]~input .bus_hold = "false";
defparam \syif.store[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N15
cycloneive_io_ibuf \syif.store[9]~input (
	.i(\syif.store [9]),
	.ibar(gnd),
	.o(\syif.store[9]~input_o ));
// synopsys translate_off
defparam \syif.store[9]~input .bus_hold = "false";
defparam \syif.store[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y0_N22
cycloneive_io_ibuf \syif.store[10]~input (
	.i(\syif.store [10]),
	.ibar(gnd),
	.o(\syif.store[10]~input_o ));
// synopsys translate_off
defparam \syif.store[10]~input .bus_hold = "false";
defparam \syif.store[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N22
cycloneive_io_ibuf \syif.store[11]~input (
	.i(\syif.store [11]),
	.ibar(gnd),
	.o(\syif.store[11]~input_o ));
// synopsys translate_off
defparam \syif.store[11]~input .bus_hold = "false";
defparam \syif.store[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y73_N1
cycloneive_io_ibuf \syif.store[12]~input (
	.i(\syif.store [12]),
	.ibar(gnd),
	.o(\syif.store[12]~input_o ));
// synopsys translate_off
defparam \syif.store[12]~input .bus_hold = "false";
defparam \syif.store[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N8
cycloneive_io_ibuf \syif.store[13]~input (
	.i(\syif.store [13]),
	.ibar(gnd),
	.o(\syif.store[13]~input_o ));
// synopsys translate_off
defparam \syif.store[13]~input .bus_hold = "false";
defparam \syif.store[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y73_N15
cycloneive_io_ibuf \syif.store[14]~input (
	.i(\syif.store [14]),
	.ibar(gnd),
	.o(\syif.store[14]~input_o ));
// synopsys translate_off
defparam \syif.store[14]~input .bus_hold = "false";
defparam \syif.store[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X56_Y0_N15
cycloneive_io_ibuf \syif.store[15]~input (
	.i(\syif.store [15]),
	.ibar(gnd),
	.o(\syif.store[15]~input_o ));
// synopsys translate_off
defparam \syif.store[15]~input .bus_hold = "false";
defparam \syif.store[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y30_N1
cycloneive_io_ibuf \syif.store[16]~input (
	.i(\syif.store [16]),
	.ibar(gnd),
	.o(\syif.store[16]~input_o ));
// synopsys translate_off
defparam \syif.store[16]~input .bus_hold = "false";
defparam \syif.store[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N15
cycloneive_io_ibuf \syif.store[17]~input (
	.i(\syif.store [17]),
	.ibar(gnd),
	.o(\syif.store[17]~input_o ));
// synopsys translate_off
defparam \syif.store[17]~input .bus_hold = "false";
defparam \syif.store[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N1
cycloneive_io_ibuf \syif.store[18]~input (
	.i(\syif.store [18]),
	.ibar(gnd),
	.o(\syif.store[18]~input_o ));
// synopsys translate_off
defparam \syif.store[18]~input .bus_hold = "false";
defparam \syif.store[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y73_N8
cycloneive_io_ibuf \syif.store[19]~input (
	.i(\syif.store [19]),
	.ibar(gnd),
	.o(\syif.store[19]~input_o ));
// synopsys translate_off
defparam \syif.store[19]~input .bus_hold = "false";
defparam \syif.store[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y73_N1
cycloneive_io_ibuf \syif.store[20]~input (
	.i(\syif.store [20]),
	.ibar(gnd),
	.o(\syif.store[20]~input_o ));
// synopsys translate_off
defparam \syif.store[20]~input .bus_hold = "false";
defparam \syif.store[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y34_N22
cycloneive_io_ibuf \syif.store[21]~input (
	.i(\syif.store [21]),
	.ibar(gnd),
	.o(\syif.store[21]~input_o ));
// synopsys translate_off
defparam \syif.store[21]~input .bus_hold = "false";
defparam \syif.store[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N22
cycloneive_io_ibuf \syif.store[22]~input (
	.i(\syif.store [22]),
	.ibar(gnd),
	.o(\syif.store[22]~input_o ));
// synopsys translate_off
defparam \syif.store[22]~input .bus_hold = "false";
defparam \syif.store[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y0_N8
cycloneive_io_ibuf \syif.store[23]~input (
	.i(\syif.store [23]),
	.ibar(gnd),
	.o(\syif.store[23]~input_o ));
// synopsys translate_off
defparam \syif.store[23]~input .bus_hold = "false";
defparam \syif.store[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y42_N15
cycloneive_io_ibuf \syif.store[24]~input (
	.i(\syif.store [24]),
	.ibar(gnd),
	.o(\syif.store[24]~input_o ));
// synopsys translate_off
defparam \syif.store[24]~input .bus_hold = "false";
defparam \syif.store[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y73_N22
cycloneive_io_ibuf \syif.store[25]~input (
	.i(\syif.store [25]),
	.ibar(gnd),
	.o(\syif.store[25]~input_o ));
// synopsys translate_off
defparam \syif.store[25]~input .bus_hold = "false";
defparam \syif.store[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X31_Y73_N8
cycloneive_io_ibuf \syif.store[26]~input (
	.i(\syif.store [26]),
	.ibar(gnd),
	.o(\syif.store[26]~input_o ));
// synopsys translate_off
defparam \syif.store[26]~input .bus_hold = "false";
defparam \syif.store[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y73_N1
cycloneive_io_ibuf \syif.store[27]~input (
	.i(\syif.store [27]),
	.ibar(gnd),
	.o(\syif.store[27]~input_o ));
// synopsys translate_off
defparam \syif.store[27]~input .bus_hold = "false";
defparam \syif.store[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N1
cycloneive_io_ibuf \syif.store[28]~input (
	.i(\syif.store [28]),
	.ibar(gnd),
	.o(\syif.store[28]~input_o ));
// synopsys translate_off
defparam \syif.store[28]~input .bus_hold = "false";
defparam \syif.store[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N15
cycloneive_io_ibuf \syif.store[29]~input (
	.i(\syif.store [29]),
	.ibar(gnd),
	.o(\syif.store[29]~input_o ));
// synopsys translate_off
defparam \syif.store[29]~input .bus_hold = "false";
defparam \syif.store[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N1
cycloneive_io_ibuf \syif.store[30]~input (
	.i(\syif.store [30]),
	.ibar(gnd),
	.o(\syif.store[30]~input_o ));
// synopsys translate_off
defparam \syif.store[30]~input .bus_hold = "false";
defparam \syif.store[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y0_N22
cycloneive_io_ibuf \syif.store[31]~input (
	.i(\syif.store [31]),
	.ibar(gnd),
	.o(\syif.store[31]~input_o ));
// synopsys translate_off
defparam \syif.store[31]~input .bus_hold = "false";
defparam \syif.store[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: CLKCTRL_G4
cycloneive_clkctrl \altera_internal_jtag~TCKUTAPclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\altera_internal_jtag~TCKUTAP }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ));
// synopsys translate_off
defparam \altera_internal_jtag~TCKUTAPclkctrl .clock_type = "global clock";
defparam \altera_internal_jtag~TCKUTAPclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G11
cycloneive_clkctrl \CPUCLK~clkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CPUCLK~q }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CPUCLK~clkctrl_outclk ));
// synopsys translate_off
defparam \CPUCLK~clkctrl .clock_type = "global clock";
defparam \CPUCLK~clkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G1
cycloneive_clkctrl \nRST~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\nRST~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\nRST~inputclkctrl_outclk ));
// synopsys translate_off
defparam \nRST~inputclkctrl .clock_type = "global clock";
defparam \nRST~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G2
cycloneive_clkctrl \CLK~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CLK~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CLK~inputclkctrl_outclk ));
// synopsys translate_off
defparam \CLK~inputclkctrl .clock_type = "global clock";
defparam \CLK~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y39_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y39_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N16
cycloneive_io_obuf \syif.halt~output (
	.i(\CPU|DP|dpif.halt~q ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.halt ),
	.obar());
// synopsys translate_off
defparam \syif.halt~output .bus_hold = "false";
defparam \syif.halt~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y0_N16
cycloneive_io_obuf \syif.load[0]~output (
	.i(\RAM|ramif.ramload[0]~0_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [0]),
	.obar());
// synopsys translate_off
defparam \syif.load[0]~output .bus_hold = "false";
defparam \syif.load[0]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X87_Y73_N16
cycloneive_io_obuf \syif.load[1]~output (
	.i(\RAM|ramif.ramload[1]~1_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [1]),
	.obar());
// synopsys translate_off
defparam \syif.load[1]~output .bus_hold = "false";
defparam \syif.load[1]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y73_N9
cycloneive_io_obuf \syif.load[2]~output (
	.i(\RAM|ramif.ramload[2]~2_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [2]),
	.obar());
// synopsys translate_off
defparam \syif.load[2]~output .bus_hold = "false";
defparam \syif.load[2]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X38_Y73_N16
cycloneive_io_obuf \syif.load[3]~output (
	.i(\RAM|ramif.ramload[3]~3_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [3]),
	.obar());
// synopsys translate_off
defparam \syif.load[3]~output .bus_hold = "false";
defparam \syif.load[3]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N16
cycloneive_io_obuf \syif.load[4]~output (
	.i(\RAM|ramif.ramload[4]~4_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [4]),
	.obar());
// synopsys translate_off
defparam \syif.load[4]~output .bus_hold = "false";
defparam \syif.load[4]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N16
cycloneive_io_obuf \syif.load[5]~output (
	.i(\RAM|ramif.ramload[5]~5_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [5]),
	.obar());
// synopsys translate_off
defparam \syif.load[5]~output .bus_hold = "false";
defparam \syif.load[5]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X72_Y73_N16
cycloneive_io_obuf \syif.load[6]~output (
	.i(\RAM|ramif.ramload[6]~6_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [6]),
	.obar());
// synopsys translate_off
defparam \syif.load[6]~output .bus_hold = "false";
defparam \syif.load[6]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y42_N2
cycloneive_io_obuf \syif.load[7]~output (
	.i(\RAM|ramif.ramload[7]~7_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [7]),
	.obar());
// synopsys translate_off
defparam \syif.load[7]~output .bus_hold = "false";
defparam \syif.load[7]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N9
cycloneive_io_obuf \syif.load[8]~output (
	.i(\RAM|ramif.ramload[8]~8_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [8]),
	.obar());
// synopsys translate_off
defparam \syif.load[8]~output .bus_hold = "false";
defparam \syif.load[8]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N2
cycloneive_io_obuf \syif.load[9]~output (
	.i(\RAM|ramif.ramload[9]~9_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [9]),
	.obar());
// synopsys translate_off
defparam \syif.load[9]~output .bus_hold = "false";
defparam \syif.load[9]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X67_Y0_N16
cycloneive_io_obuf \syif.load[10]~output (
	.i(\RAM|ramif.ramload[10]~10_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [10]),
	.obar());
// synopsys translate_off
defparam \syif.load[10]~output .bus_hold = "false";
defparam \syif.load[10]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N9
cycloneive_io_obuf \syif.load[11]~output (
	.i(\RAM|ramif.ramload[11]~11_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [11]),
	.obar());
// synopsys translate_off
defparam \syif.load[11]~output .bus_hold = "false";
defparam \syif.load[11]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N23
cycloneive_io_obuf \syif.load[12]~output (
	.i(\RAM|ramif.ramload[12]~12_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [12]),
	.obar());
// synopsys translate_off
defparam \syif.load[12]~output .bus_hold = "false";
defparam \syif.load[12]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X67_Y73_N23
cycloneive_io_obuf \syif.load[13]~output (
	.i(\RAM|ramif.ramload[13]~13_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [13]),
	.obar());
// synopsys translate_off
defparam \syif.load[13]~output .bus_hold = "false";
defparam \syif.load[13]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X38_Y73_N23
cycloneive_io_obuf \syif.load[14]~output (
	.i(\RAM|ramif.ramload[14]~14_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [14]),
	.obar());
// synopsys translate_off
defparam \syif.load[14]~output .bus_hold = "false";
defparam \syif.load[14]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X72_Y73_N9
cycloneive_io_obuf \syif.load[15]~output (
	.i(\RAM|ramif.ramload[15]~15_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [15]),
	.obar());
// synopsys translate_off
defparam \syif.load[15]~output .bus_hold = "false";
defparam \syif.load[15]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y0_N23
cycloneive_io_obuf \syif.load[16]~output (
	.i(\RAM|ramif.ramload[16]~17_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [16]),
	.obar());
// synopsys translate_off
defparam \syif.load[16]~output .bus_hold = "false";
defparam \syif.load[16]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y33_N2
cycloneive_io_obuf \syif.load[17]~output (
	.i(\RAM|ramif.ramload[17]~19_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [17]),
	.obar());
// synopsys translate_off
defparam \syif.load[17]~output .bus_hold = "false";
defparam \syif.load[17]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y0_N2
cycloneive_io_obuf \syif.load[18]~output (
	.i(\RAM|ramif.ramload[18]~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [18]),
	.obar());
// synopsys translate_off
defparam \syif.load[18]~output .bus_hold = "false";
defparam \syif.load[18]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y73_N2
cycloneive_io_obuf \syif.load[19]~output (
	.i(\RAM|ramif.ramload[19]~21_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [19]),
	.obar());
// synopsys translate_off
defparam \syif.load[19]~output .bus_hold = "false";
defparam \syif.load[19]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N2
cycloneive_io_obuf \syif.load[20]~output (
	.i(\RAM|ramif.ramload[20]~22_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [20]),
	.obar());
// synopsys translate_off
defparam \syif.load[20]~output .bus_hold = "false";
defparam \syif.load[20]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y40_N9
cycloneive_io_obuf \syif.load[21]~output (
	.i(\RAM|ramif.ramload[21]~23_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [21]),
	.obar());
// synopsys translate_off
defparam \syif.load[21]~output .bus_hold = "false";
defparam \syif.load[21]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y35_N16
cycloneive_io_obuf \syif.load[22]~output (
	.i(\RAM|ramif.ramload[22]~24_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [22]),
	.obar());
// synopsys translate_off
defparam \syif.load[22]~output .bus_hold = "false";
defparam \syif.load[22]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y0_N2
cycloneive_io_obuf \syif.load[23]~output (
	.i(\RAM|ramif.ramload[23]~25_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [23]),
	.obar());
// synopsys translate_off
defparam \syif.load[23]~output .bus_hold = "false";
defparam \syif.load[23]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y34_N23
cycloneive_io_obuf \syif.load[24]~output (
	.i(\RAM|ramif.ramload[24]~26_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [24]),
	.obar());
// synopsys translate_off
defparam \syif.load[24]~output .bus_hold = "false";
defparam \syif.load[24]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X47_Y0_N2
cycloneive_io_obuf \syif.load[25]~output (
	.i(\RAM|ramif.ramload[25]~27_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [25]),
	.obar());
// synopsys translate_off
defparam \syif.load[25]~output .bus_hold = "false";
defparam \syif.load[25]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N23
cycloneive_io_obuf \syif.load[26]~output (
	.i(\RAM|ramif.ramload[26]~28_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [26]),
	.obar());
// synopsys translate_off
defparam \syif.load[26]~output .bus_hold = "false";
defparam \syif.load[26]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y0_N9
cycloneive_io_obuf \syif.load[27]~output (
	.i(\RAM|ramif.ramload[27]~29_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [27]),
	.obar());
// synopsys translate_off
defparam \syif.load[27]~output .bus_hold = "false";
defparam \syif.load[27]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X40_Y73_N9
cycloneive_io_obuf \syif.load[28]~output (
	.i(\RAM|ramif.ramload[28]~30_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [28]),
	.obar());
// synopsys translate_off
defparam \syif.load[28]~output .bus_hold = "false";
defparam \syif.load[28]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y0_N2
cycloneive_io_obuf \syif.load[29]~output (
	.i(\RAM|ramif.ramload[29]~31_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [29]),
	.obar());
// synopsys translate_off
defparam \syif.load[29]~output .bus_hold = "false";
defparam \syif.load[29]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N9
cycloneive_io_obuf \syif.load[30]~output (
	.i(\RAM|ramif.ramload[30]~32_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [30]),
	.obar());
// synopsys translate_off
defparam \syif.load[30]~output .bus_hold = "false";
defparam \syif.load[30]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y0_N16
cycloneive_io_obuf \syif.load[31]~output (
	.i(\RAM|ramif.ramload[31]~33_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [31]),
	.obar());
// synopsys translate_off
defparam \syif.load[31]~output .bus_hold = "false";
defparam \syif.load[31]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y37_N1
cycloneive_io_obuf \altera_reserved_tdo~output (
	.i(\altera_internal_jtag~TDO ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(altera_reserved_tdo),
	.obar());
// synopsys translate_off
defparam \altera_reserved_tdo~output .bus_hold = "false";
defparam \altera_reserved_tdo~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOIBUF_X0_Y38_N1
cycloneive_io_ibuf \altera_reserved_tms~input (
	.i(altera_reserved_tms),
	.ibar(gnd),
	.o(\altera_reserved_tms~input_o ));
// synopsys translate_off
defparam \altera_reserved_tms~input .bus_hold = "false";
defparam \altera_reserved_tms~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y39_N1
cycloneive_io_ibuf \altera_reserved_tck~input (
	.i(altera_reserved_tck),
	.ibar(gnd),
	.o(\altera_reserved_tck~input_o ));
// synopsys translate_off
defparam \altera_reserved_tck~input .bus_hold = "false";
defparam \altera_reserved_tck~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y40_N1
cycloneive_io_ibuf \altera_reserved_tdi~input (
	.i(altera_reserved_tdi),
	.ibar(gnd),
	.o(\altera_reserved_tdi~input_o ));
// synopsys translate_off
defparam \altera_reserved_tdi~input .bus_hold = "false";
defparam \altera_reserved_tdi~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 .lut_mask = 16'h33CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~10 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9 .lut_mask = 16'hC303;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13 .lut_mask = 16'hC303;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .lut_mask = 16'hCC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y41_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .lut_mask = 16'hFA00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hF0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .lut_mask = 16'hF0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .lut_mask = 16'hF0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .lut_mask = 16'hF0E0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y40_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y41_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .lut_mask = 16'h0A0A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y41_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y41_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y41_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y41_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .lut_mask = 16'h3CF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y41_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .lut_mask = 16'h5575;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .lut_mask = 16'hFEFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y40_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y40_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y40_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y40_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y40_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .lut_mask = 16'h0001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y40_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y40_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y40_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y40_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y40_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y40_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y40_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y40_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y40_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y40_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y40_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y40_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y40_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y40_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y40_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .lut_mask = 16'h0008;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y40_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y40_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8 .lut_mask = 16'hF888;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y39_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 .lut_mask = 16'h5A5A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X36_Y39_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X35_Y39_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .lut_mask = 16'h0003;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y39_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .lut_mask = 16'hCC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7 .lut_mask = 16'hFF04;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y39_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X36_Y39_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~7_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12 .lut_mask = 16'h8000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X35_Y39_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .lut_mask = 16'h0197;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y39_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 .lut_mask = 16'hCC48;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y39_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .lut_mask = 16'hBB88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y39_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .lut_mask = 16'hFFFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(gnd),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .lut_mask = 16'hD8D8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N22
cycloneive_lcell_comb \~QIC_CREATED_GND~I (
// Equation(s):
// \~QIC_CREATED_GND~I_combout  = GND

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~QIC_CREATED_GND~I_combout ),
	.cout());
// synopsys translate_off
defparam \~QIC_CREATED_GND~I .lut_mask = 16'h0000;
defparam \~QIC_CREATED_GND~I .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y41_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.asdata(\~QIC_CREATED_GND~I_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .lut_mask = 16'hFC30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .lut_mask = 16'hC080;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .lut_mask = 16'h30B8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y41_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y41_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.datac(gnd),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .lut_mask = 16'hEE44;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .lut_mask = 16'hFC30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y41_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y41_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .lut_mask = 16'hF3C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y41_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .lut_mask = 16'hFC0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .lut_mask = 16'hC840;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y41_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .lut_mask = 16'h41C8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .lut_mask = 16'hD2F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y41_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y41_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .lut_mask = 16'h2000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y39_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .lut_mask = 16'h50D8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y39_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y41_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .lut_mask = 16'hFFFD;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y41_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y39_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y39_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y41_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .lut_mask = 16'hFC30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y41_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y40_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .lut_mask = 16'h0800;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y39_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .lut_mask = 16'h00C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y39_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y39_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y39_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y39_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y39_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y39_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y39_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .lut_mask = 16'h0008;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y39_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y39_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y39_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y39_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y39_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y39_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y39_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y39_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y40_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .lut_mask = 16'h0800;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y40_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y39_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .lut_mask = 16'h3F3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y39_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .lut_mask = 16'hFC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y39_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X39_Y39_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X39_Y39_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X39_Y39_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y40_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .lut_mask = 16'h00F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y40_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y40_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y40_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .lut_mask = 16'hFFCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y40_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y40_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .lut_mask = 16'h3030;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y40_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y40_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .lut_mask = 16'hFFCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y40_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h33CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .lut_mask = 16'hC30C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h3C3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .lut_mask = 16'hFF40;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y40_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .lut_mask = 16'hA5A5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X41_Y40_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .lut_mask = 16'hFFFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .lut_mask = 16'hAE0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y40_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .lut_mask = 16'h3C3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X41_Y40_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y40_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .lut_mask = 16'hA3A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .lut_mask = 16'h44CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .lut_mask = 16'hFFC8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y40_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .lut_mask = 16'hA001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .lut_mask = 16'h0004;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .lut_mask = 16'hF0F8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y40_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y40_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .lut_mask = 16'hADA8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y39_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .lut_mask = 16'hFC30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y39_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y40_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .lut_mask = 16'hAAE4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y40_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .lut_mask = 16'h1A5F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y40_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo (
	.clk(!\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X16_Y38_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y66_N0
cycloneive_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y40_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y40_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module ram (
	is_in_use_reg,
	ramaddr,
	ramaddr1,
	ramaddr2,
	ramaddr3,
	ramaddr4,
	ramaddr5,
	ramaddr6,
	ramaddr7,
	ramaddr8,
	ramaddr9,
	ramaddr10,
	ramaddr11,
	ramaddr12,
	ramaddr13,
	ramaddr14,
	ramaddr15,
	\ramif.ramaddr ,
	ramaddr16,
	ramaddr17,
	ramaddr18,
	ramaddr19,
	ramaddr20,
	ramaddr21,
	ramaddr22,
	ramaddr23,
	ramaddr24,
	\ramif.ramWEN ,
	\ramif.ramREN ,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	ramstore,
	ramstore1,
	ramstore2,
	ramstore3,
	ramstore4,
	ramstore5,
	ramstore6,
	ramstore7,
	ramstore8,
	ramstore9,
	ramstore10,
	ramstore11,
	ramstore12,
	ramstore13,
	ramstore14,
	ramstore15,
	ramstore16,
	ramstore17,
	ramstore18,
	ramstore19,
	ramstore20,
	ramstore21,
	ramstore22,
	ramstore23,
	ramstore24,
	ramstore25,
	ramstore26,
	ramstore27,
	ramstore28,
	ramstore29,
	ramstore30,
	ramstore31,
	ramaddr25,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	nRST,
	altera_internal_jtag1,
	nRST1,
	CLK,
	devpor,
	devclrn,
	devoe);
output 	is_in_use_reg;
input 	ramaddr;
input 	ramaddr1;
input 	ramaddr2;
input 	ramaddr3;
input 	ramaddr4;
input 	ramaddr5;
input 	ramaddr6;
input 	ramaddr7;
input 	ramaddr8;
input 	ramaddr9;
input 	ramaddr10;
input 	ramaddr11;
input 	ramaddr12;
input 	ramaddr13;
input 	ramaddr14;
input 	ramaddr15;
input 	[31:0] \ramif.ramaddr ;
input 	ramaddr16;
input 	ramaddr17;
input 	ramaddr18;
input 	ramaddr19;
input 	ramaddr20;
input 	ramaddr21;
input 	ramaddr22;
input 	ramaddr23;
input 	ramaddr24;
input 	\ramif.ramWEN ;
input 	\ramif.ramREN ;
output 	always1;
output 	ramiframload_0;
output 	ramiframload_1;
output 	ramiframload_2;
output 	ramiframload_3;
output 	ramiframload_4;
output 	ramiframload_5;
output 	ramiframload_6;
output 	ramiframload_7;
output 	ramiframload_8;
output 	ramiframload_9;
output 	ramiframload_10;
output 	ramiframload_11;
output 	ramiframload_12;
output 	ramiframload_13;
output 	ramiframload_14;
output 	ramiframload_15;
output 	ramiframload_16;
output 	ramiframload_17;
output 	ramiframload_18;
output 	ramiframload_19;
output 	ramiframload_20;
output 	ramiframload_21;
output 	ramiframload_22;
output 	ramiframload_23;
output 	ramiframload_24;
output 	ramiframload_25;
output 	ramiframload_26;
output 	ramiframload_27;
output 	ramiframload_28;
output 	ramiframload_29;
output 	ramiframload_30;
output 	ramiframload_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	ramstore;
input 	ramstore1;
input 	ramstore2;
input 	ramstore3;
input 	ramstore4;
input 	ramstore5;
input 	ramstore6;
input 	ramstore7;
input 	ramstore8;
input 	ramstore9;
input 	ramstore10;
input 	ramstore11;
input 	ramstore12;
input 	ramstore13;
input 	ramstore14;
input 	ramstore15;
input 	ramstore16;
input 	ramstore17;
input 	ramstore18;
input 	ramstore19;
input 	ramstore20;
input 	ramstore21;
input 	ramstore22;
input 	ramstore23;
input 	ramstore24;
input 	ramstore25;
input 	ramstore26;
input 	ramstore27;
input 	ramstore28;
input 	ramstore29;
input 	ramstore30;
input 	ramstore31;
input 	ramaddr25;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	nRST;
input 	altera_internal_jtag1;
input 	nRST1;
input 	CLK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ;
wire \Equal2~1_combout ;
wire \Equal2~7_combout ;
wire \Equal2~10_combout ;
wire \Equal2~15_combout ;
wire \always0~0_combout ;
wire \addr[7]~feeder_combout ;
wire \addr[11]~feeder_combout ;
wire \always0~1_combout ;
wire \Equal2~18_combout ;
wire \Equal2~16_combout ;
wire \Equal2~17_combout ;
wire \Equal2~19_combout ;
wire \Equal2~11_combout ;
wire \Equal2~13_combout ;
wire \Equal2~12_combout ;
wire \Equal2~14_combout ;
wire \Equal2~6_combout ;
wire \Equal2~5_combout ;
wire \Equal2~8_combout ;
wire \Equal2~9_combout ;
wire \Equal2~2_combout ;
wire \Equal2~0_combout ;
wire \Equal2~3_combout ;
wire \Equal2~4_combout ;
wire \Equal2~20_combout ;
wire \ramif.ramload[16]~16_combout ;
wire \ramif.ramload[17]~18_combout ;
wire [1:0] en;
wire [31:0] addr;
wire [0:0] \altsyncram_component|auto_generated|altsyncram1|address_reg_a ;


altsyncram_1 altsyncram_component(
	.ram_block3a32(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.ram_block3a0(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.ram_block3a33(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.ram_block3a1(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.ram_block3a34(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.ram_block3a2(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.ram_block3a35(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.ram_block3a3(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.ram_block3a36(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.ram_block3a4(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.ram_block3a37(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.ram_block3a5(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.ram_block3a38(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.ram_block3a6(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.ram_block3a39(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.ram_block3a7(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.ram_block3a40(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.ram_block3a8(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.ram_block3a41(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.ram_block3a9(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.ram_block3a42(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.ram_block3a10(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.ram_block3a43(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.ram_block3a11(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.ram_block3a44(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.ram_block3a12(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.ram_block3a45(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.ram_block3a13(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.ram_block3a46(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.ram_block3a14(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.ram_block3a47(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.ram_block3a15(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.ram_block3a48(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.ram_block3a16(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.ram_block3a49(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.ram_block3a17(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.ram_block3a50(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.ram_block3a18(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.ram_block3a51(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.ram_block3a19(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.ram_block3a52(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.ram_block3a20(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.ram_block3a53(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.ram_block3a21(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.ram_block3a54(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.ram_block3a22(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.ram_block3a55(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.ram_block3a23(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.ram_block3a56(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.ram_block3a24(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.ram_block3a57(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.ram_block3a25(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.ram_block3a58(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.ram_block3a26(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.ram_block3a59(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.ram_block3a27(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.ram_block3a60(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.ram_block3a28(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.ram_block3a61(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.ram_block3a29(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.ram_block3a62(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.ram_block3a30(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.ram_block3a63(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.ram_block3a31(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.address_a({gnd,ramaddr15,ramaddr12,ramaddr13,ramaddr10,ramaddr11,ramaddr8,ramaddr9,ramaddr6,ramaddr7,ramaddr4,ramaddr5,ramaddr2,ramaddr3}),
	.ramaddr(ramaddr14),
	.ramWEN(\ramif.ramWEN ),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.data_a({ramstore31,ramstore30,ramstore29,ramstore28,ramstore27,ramstore26,ramstore25,ramstore24,ramstore23,ramstore22,ramstore21,ramstore20,ramstore19,ramstore18,ramstore17,ramstore16,ramstore15,ramstore14,ramstore13,ramstore12,ramstore11,ramstore10,ramstore9,ramstore8,ramstore7,ramstore6,
ramstore5,ramstore4,ramstore3,ramstore2,ramstore1,ramstore}),
	.ramaddr1(ramaddr25),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(CLK),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: FF_X59_Y31_N17
dffeas \addr[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr3),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[2]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[2] .is_wysiwyg = "true";
defparam \addr[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N7
dffeas \addr[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr2),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[3]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[3] .is_wysiwyg = "true";
defparam \addr[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N16
cycloneive_lcell_comb \Equal2~1 (
// Equation(s):
// \Equal2~1_combout  = (\ramaddr~5_combout  & (addr[3] & (addr[2] $ (!\ramaddr~7_combout )))) # (!\ramaddr~5_combout  & (!addr[3] & (addr[2] $ (!\ramaddr~7_combout ))))

	.dataa(ramaddr2),
	.datab(addr[3]),
	.datac(addr[2]),
	.datad(ramaddr3),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~1 .lut_mask = 16'h9009;
defparam \Equal2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N23
dffeas \addr[5] (
	.clk(CLK),
	.d(ramaddr4),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[5]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[5] .is_wysiwyg = "true";
defparam \addr[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N7
dffeas \addr[7] (
	.clk(CLK),
	.d(\addr[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[7]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[7] .is_wysiwyg = "true";
defparam \addr[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N27
dffeas \addr[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr8),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[9]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[9] .is_wysiwyg = "true";
defparam \addr[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N23
dffeas \addr[11] (
	.clk(CLK),
	.d(\addr[11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[11]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[11] .is_wysiwyg = "true";
defparam \addr[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y35_N9
dffeas \addr[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr13),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[12]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[12] .is_wysiwyg = "true";
defparam \addr[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y35_N11
dffeas \addr[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr12),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[13]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[13] .is_wysiwyg = "true";
defparam \addr[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N8
cycloneive_lcell_comb \Equal2~7 (
// Equation(s):
// \Equal2~7_combout  = (addr[13] & (\ramaddr~25_combout  & (\ramaddr~27_combout  $ (!addr[12])))) # (!addr[13] & (!\ramaddr~25_combout  & (\ramaddr~27_combout  $ (!addr[12]))))

	.dataa(addr[13]),
	.datab(ramaddr13),
	.datac(addr[12]),
	.datad(ramaddr12),
	.cin(gnd),
	.combout(\Equal2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~7 .lut_mask = 16'h8241;
defparam \Equal2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N27
dffeas \addr[15] (
	.clk(CLK),
	.d(ramaddr25),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[15]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[15] .is_wysiwyg = "true";
defparam \addr[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y34_N15
dffeas \addr[16] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr16),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[16]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[16] .is_wysiwyg = "true";
defparam \addr[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y34_N21
dffeas \addr[17] (
	.clk(CLK),
	.d(\ramif.ramaddr [17]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[17]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[17] .is_wysiwyg = "true";
defparam \addr[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N14
cycloneive_lcell_comb \Equal2~10 (
// Equation(s):
// \Equal2~10_combout  = (addr[17] & (\ramaddr~33_combout  & (\ramaddr~35_combout  $ (!addr[16])))) # (!addr[17] & (!\ramaddr~33_combout  & (\ramaddr~35_combout  $ (!addr[16]))))

	.dataa(addr[17]),
	.datab(ramaddr16),
	.datac(addr[16]),
	.datad(\ramif.ramaddr [17]),
	.cin(gnd),
	.combout(\Equal2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~10 .lut_mask = 16'h8241;
defparam \Equal2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N19
dffeas \addr[23] (
	.clk(CLK),
	.d(\ramif.ramaddr [23]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[23]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[23] .is_wysiwyg = "true";
defparam \addr[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N13
dffeas \addr[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr21),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[24]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[24] .is_wysiwyg = "true";
defparam \addr[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N15
dffeas \addr[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr20),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[25]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[25] .is_wysiwyg = "true";
defparam \addr[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N12
cycloneive_lcell_comb \Equal2~15 (
// Equation(s):
// \Equal2~15_combout  = (\ramaddr~51_combout  & (addr[24] & (addr[25] $ (!\ramaddr~49_combout )))) # (!\ramaddr~51_combout  & (!addr[24] & (addr[25] $ (!\ramaddr~49_combout ))))

	.dataa(ramaddr21),
	.datab(addr[25]),
	.datac(addr[24]),
	.datad(ramaddr20),
	.cin(gnd),
	.combout(\Equal2~15_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~15 .lut_mask = 16'h8421;
defparam \Equal2~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N1
dffeas \en[1] (
	.clk(CLK),
	.d(\ramif.ramREN ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[1]),
	.prn(vcc));
// synopsys translate_off
defparam \en[1] .is_wysiwyg = "true";
defparam \en[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N31
dffeas \en[0] (
	.clk(CLK),
	.d(\ramif.ramWEN ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[0]),
	.prn(vcc));
// synopsys translate_off
defparam \en[0] .is_wysiwyg = "true";
defparam \en[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N10
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// \always0~0_combout  = (\ramWEN~0_combout  & ((en[1] $ (\ramREN~0_combout )) # (!en[0]))) # (!\ramWEN~0_combout  & ((en[0]) # (en[1] $ (\ramREN~0_combout ))))

	.dataa(\ramif.ramWEN ),
	.datab(en[0]),
	.datac(en[1]),
	.datad(\ramif.ramREN ),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'h6FF6;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N6
cycloneive_lcell_comb \addr[7]~feeder (
// Equation(s):
// \addr[7]~feeder_combout  = \ramaddr~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr6),
	.cin(gnd),
	.combout(\addr[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[7]~feeder .lut_mask = 16'hFF00;
defparam \addr[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N22
cycloneive_lcell_comb \addr[11]~feeder (
// Equation(s):
// \addr[11]~feeder_combout  = \ramaddr~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr10),
	.cin(gnd),
	.combout(\addr[11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[11]~feeder .lut_mask = 16'hFF00;
defparam \addr[11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N2
cycloneive_lcell_comb \always1~0 (
// Equation(s):
// always1 = ((\Equal2~20_combout  & ((!\ramREN~0_combout ) # (!\ramWEN~0_combout )))) # (!\nRST~input_o )

	.dataa(\ramif.ramWEN ),
	.datab(\ramif.ramREN ),
	.datac(nRST),
	.datad(\Equal2~20_combout ),
	.cin(gnd),
	.combout(always1),
	.cout());
// synopsys translate_off
defparam \always1~0 .lut_mask = 16'h7F0F;
defparam \always1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N22
cycloneive_lcell_comb \ramif.ramload[0]~0 (
// Equation(s):
// ramiframload_0 = ((address_reg_a_0 & (ram_block3a321)) # (!address_reg_a_0 & ((ram_block3a01)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.cin(gnd),
	.combout(ramiframload_0),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[0]~0 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N8
cycloneive_lcell_comb \ramif.ramload[1]~1 (
// Equation(s):
// ramiframload_1 = (always1 & ((address_reg_a_0 & (ram_block3a331)) # (!address_reg_a_0 & ((ram_block3a110)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.cin(gnd),
	.combout(ramiframload_1),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[1]~1 .lut_mask = 16'hC480;
defparam \ramif.ramload[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N12
cycloneive_lcell_comb \ramif.ramload[2]~2 (
// Equation(s):
// ramiframload_2 = (always1 & ((address_reg_a_0 & (ram_block3a341)) # (!address_reg_a_0 & ((ram_block3a210)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_2),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[2]~2 .lut_mask = 16'hD800;
defparam \ramif.ramload[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N14
cycloneive_lcell_comb \ramif.ramload[3]~3 (
// Equation(s):
// ramiframload_3 = (always1 & ((address_reg_a_0 & (ram_block3a351)) # (!address_reg_a_0 & ((ram_block3a310)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_3),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[3]~3 .lut_mask = 16'hAC00;
defparam \ramif.ramload[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N12
cycloneive_lcell_comb \ramif.ramload[4]~4 (
// Equation(s):
// ramiframload_4 = ((address_reg_a_0 & ((ram_block3a361))) # (!address_reg_a_0 & (ram_block3a410))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.cin(gnd),
	.combout(ramiframload_4),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[4]~4 .lut_mask = 16'hFD5D;
defparam \ramif.ramload[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N14
cycloneive_lcell_comb \ramif.ramload[5]~5 (
// Equation(s):
// ramiframload_5 = (always1 & ((address_reg_a_0 & (ram_block3a371)) # (!address_reg_a_0 & ((ram_block3a510)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.cin(gnd),
	.combout(ramiframload_5),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[5]~5 .lut_mask = 16'hD080;
defparam \ramif.ramload[5]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N0
cycloneive_lcell_comb \ramif.ramload[6]~6 (
// Equation(s):
// ramiframload_6 = ((address_reg_a_0 & (ram_block3a381)) # (!address_reg_a_0 & ((ram_block3a64)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.cin(gnd),
	.combout(ramiframload_6),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[6]~6 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[6]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N22
cycloneive_lcell_comb \ramif.ramload[7]~7 (
// Equation(s):
// ramiframload_7 = ((address_reg_a_0 & ((ram_block3a391))) # (!address_reg_a_0 & (ram_block3a71))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.cin(gnd),
	.combout(ramiframload_7),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[7]~7 .lut_mask = 16'hFD75;
defparam \ramif.ramload[7]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N30
cycloneive_lcell_comb \ramif.ramload[8]~8 (
// Equation(s):
// ramiframload_8 = (always1 & ((address_reg_a_0 & ((ram_block3a401))) # (!address_reg_a_0 & (ram_block3a81))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.cin(gnd),
	.combout(ramiframload_8),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[8]~8 .lut_mask = 16'hE020;
defparam \ramif.ramload[8]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N28
cycloneive_lcell_comb \ramif.ramload[9]~9 (
// Equation(s):
// ramiframload_9 = ((address_reg_a_0 & ((ram_block3a412))) # (!address_reg_a_0 & (ram_block3a91))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.cin(gnd),
	.combout(ramiframload_9),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[9]~9 .lut_mask = 16'hFD75;
defparam \ramif.ramload[9]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N26
cycloneive_lcell_comb \ramif.ramload[10]~10 (
// Equation(s):
// ramiframload_10 = (always1 & ((address_reg_a_0 & ((ram_block3a421))) # (!address_reg_a_0 & (ram_block3a101))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.cin(gnd),
	.combout(ramiframload_10),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[10]~10 .lut_mask = 16'hE020;
defparam \ramif.ramload[10]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N10
cycloneive_lcell_comb \ramif.ramload[11]~11 (
// Equation(s):
// ramiframload_11 = ((address_reg_a_0 & (ram_block3a431)) # (!address_reg_a_0 & ((ram_block3a112)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.cin(gnd),
	.combout(ramiframload_11),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[11]~11 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[11]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N0
cycloneive_lcell_comb \ramif.ramload[12]~12 (
// Equation(s):
// ramiframload_12 = ((address_reg_a_0 & (ram_block3a441)) # (!address_reg_a_0 & ((ram_block3a121)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.cin(gnd),
	.combout(ramiframload_12),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[12]~12 .lut_mask = 16'hF7D5;
defparam \ramif.ramload[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N12
cycloneive_lcell_comb \ramif.ramload[13]~13 (
// Equation(s):
// ramiframload_13 = ((address_reg_a_0 & ((ram_block3a451))) # (!address_reg_a_0 & (ram_block3a131))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.cin(gnd),
	.combout(ramiframload_13),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[13]~13 .lut_mask = 16'hFB73;
defparam \ramif.ramload[13]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N18
cycloneive_lcell_comb \ramif.ramload[14]~14 (
// Equation(s):
// ramiframload_14 = (always1 & ((address_reg_a_0 & (ram_block3a461)) # (!address_reg_a_0 & ((ram_block3a141)))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.cin(gnd),
	.combout(ramiframload_14),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[14]~14 .lut_mask = 16'h8A80;
defparam \ramif.ramload[14]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N2
cycloneive_lcell_comb \ramif.ramload[15]~15 (
// Equation(s):
// ramiframload_15 = ((address_reg_a_0 & ((ram_block3a471))) # (!address_reg_a_0 & (ram_block3a151))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.cin(gnd),
	.combout(ramiframload_15),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[15]~15 .lut_mask = 16'hFB73;
defparam \ramif.ramload[15]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N4
cycloneive_lcell_comb \ramif.ramload[16]~17 (
// Equation(s):
// ramiframload_16 = (\ramif.ramload[16]~16_combout ) # ((address_reg_a_0 & ((ram_block3a481))) # (!address_reg_a_0 & (ram_block3a161)))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.datab(\ramif.ramload[16]~16_combout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.cin(gnd),
	.combout(ramiframload_16),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[16]~17 .lut_mask = 16'hFECE;
defparam \ramif.ramload[16]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N24
cycloneive_lcell_comb \ramif.ramload[17]~19 (
// Equation(s):
// ramiframload_17 = (!\ramif.ramload[17]~18_combout  & ((address_reg_a_0 & ((ram_block3a491))) # (!address_reg_a_0 & (ram_block3a171))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\ramif.ramload[17]~18_combout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.cin(gnd),
	.combout(ramiframload_17),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[17]~19 .lut_mask = 16'h0E02;
defparam \ramif.ramload[17]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N10
cycloneive_lcell_comb \ramif.ramload[18]~20 (
// Equation(s):
// ramiframload_18 = (always1 & ((address_reg_a_0 & ((ram_block3a501))) # (!address_reg_a_0 & (ram_block3a181))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.cin(gnd),
	.combout(ramiframload_18),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[18]~20 .lut_mask = 16'hA820;
defparam \ramif.ramload[18]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N30
cycloneive_lcell_comb \ramif.ramload[19]~21 (
// Equation(s):
// ramiframload_19 = (always1 & ((address_reg_a_0 & (ram_block3a512)) # (!address_reg_a_0 & ((ram_block3a191)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.cin(gnd),
	.combout(ramiframload_19),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[19]~21 .lut_mask = 16'hD080;
defparam \ramif.ramload[19]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N8
cycloneive_lcell_comb \ramif.ramload[20]~22 (
// Equation(s):
// ramiframload_20 = ((address_reg_a_0 & (ram_block3a521)) # (!address_reg_a_0 & ((ram_block3a201)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.cin(gnd),
	.combout(ramiframload_20),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[20]~22 .lut_mask = 16'hBF8F;
defparam \ramif.ramload[20]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N6
cycloneive_lcell_comb \ramif.ramload[21]~23 (
// Equation(s):
// ramiframload_21 = (always1 & ((address_reg_a_0 & ((ram_block3a531))) # (!address_reg_a_0 & (ram_block3a212))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_21),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[21]~23 .lut_mask = 16'hE400;
defparam \ramif.ramload[21]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N18
cycloneive_lcell_comb \ramif.ramload[22]~24 (
// Equation(s):
// ramiframload_22 = ((address_reg_a_0 & ((ram_block3a541))) # (!address_reg_a_0 & (ram_block3a221))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.cin(gnd),
	.combout(ramiframload_22),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[22]~24 .lut_mask = 16'hEF4F;
defparam \ramif.ramload[22]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N10
cycloneive_lcell_comb \ramif.ramload[23]~25 (
// Equation(s):
// ramiframload_23 = ((address_reg_a_0 & ((ram_block3a551))) # (!address_reg_a_0 & (ram_block3a231))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.cin(gnd),
	.combout(ramiframload_23),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[23]~25 .lut_mask = 16'hFB73;
defparam \ramif.ramload[23]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N28
cycloneive_lcell_comb \ramif.ramload[24]~26 (
// Equation(s):
// ramiframload_24 = (always1 & ((address_reg_a_0 & ((ram_block3a561))) # (!address_reg_a_0 & (ram_block3a241))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.cin(gnd),
	.combout(ramiframload_24),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[24]~26 .lut_mask = 16'hC840;
defparam \ramif.ramload[24]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N8
cycloneive_lcell_comb \ramif.ramload[25]~27 (
// Equation(s):
// ramiframload_25 = ((address_reg_a_0 & ((ram_block3a571))) # (!address_reg_a_0 & (ram_block3a251))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.cin(gnd),
	.combout(ramiframload_25),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[25]~27 .lut_mask = 16'hEF4F;
defparam \ramif.ramload[25]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N20
cycloneive_lcell_comb \ramif.ramload[26]~28 (
// Equation(s):
// ramiframload_26 = (always1 & ((address_reg_a_0 & (ram_block3a581)) # (!address_reg_a_0 & ((ram_block3a261)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_26),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[26]~28 .lut_mask = 16'hD800;
defparam \ramif.ramload[26]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N6
cycloneive_lcell_comb \ramif.ramload[27]~29 (
// Equation(s):
// ramiframload_27 = ((address_reg_a_0 & (ram_block3a591)) # (!address_reg_a_0 & ((ram_block3a271)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.cin(gnd),
	.combout(ramiframload_27),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[27]~29 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[27]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N14
cycloneive_lcell_comb \ramif.ramload[28]~30 (
// Equation(s):
// ramiframload_28 = ((address_reg_a_0 & (ram_block3a601)) # (!address_reg_a_0 & ((ram_block3a281)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_28),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[28]~30 .lut_mask = 16'hD8FF;
defparam \ramif.ramload[28]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N12
cycloneive_lcell_comb \ramif.ramload[29]~31 (
// Equation(s):
// ramiframload_29 = (\ramif.ramload[16]~16_combout ) # ((address_reg_a_0 & (ram_block3a611)) # (!address_reg_a_0 & ((ram_block3a291))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\ramif.ramload[16]~16_combout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.cin(gnd),
	.combout(ramiframload_29),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[29]~31 .lut_mask = 16'hFDEC;
defparam \ramif.ramload[29]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N8
cycloneive_lcell_comb \ramif.ramload[30]~32 (
// Equation(s):
// ramiframload_30 = (always1 & ((address_reg_a_0 & (ram_block3a621)) # (!address_reg_a_0 & ((ram_block3a301)))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.cin(gnd),
	.combout(ramiframload_30),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[30]~32 .lut_mask = 16'hA280;
defparam \ramif.ramload[30]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N2
cycloneive_lcell_comb \ramif.ramload[31]~33 (
// Equation(s):
// ramiframload_31 = ((address_reg_a_0 & (ram_block3a631)) # (!address_reg_a_0 & ((ram_block3a312)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.cin(gnd),
	.combout(ramiframload_31),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[31]~33 .lut_mask = 16'hF7D5;
defparam \ramif.ramload[31]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N22
cycloneive_lcell_comb \always0~1 (
// Equation(s):
// \always0~1_combout  = (\always0~0_combout ) # (((\ramREN~0_combout  & \ramWEN~0_combout )) # (!\Equal2~20_combout ))

	.dataa(\always0~0_combout ),
	.datab(\ramif.ramREN ),
	.datac(\ramif.ramWEN ),
	.datad(\Equal2~20_combout ),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
// synopsys translate_off
defparam \always0~1 .lut_mask = 16'hEAFF;
defparam \always0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N29
dffeas \addr[30] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr24),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[30]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[30] .is_wysiwyg = "true";
defparam \addr[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N15
dffeas \addr[31] (
	.clk(CLK),
	.d(\ramif.ramaddr [31]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[31]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[31] .is_wysiwyg = "true";
defparam \addr[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N28
cycloneive_lcell_comb \Equal2~18 (
// Equation(s):
// \Equal2~18_combout  = (\ramaddr~63_combout  & (addr[30] & (\ramaddr~61_combout  $ (!addr[31])))) # (!\ramaddr~63_combout  & (!addr[30] & (\ramaddr~61_combout  $ (!addr[31]))))

	.dataa(ramaddr24),
	.datab(\ramif.ramaddr [31]),
	.datac(addr[30]),
	.datad(addr[31]),
	.cin(gnd),
	.combout(\Equal2~18_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~18 .lut_mask = 16'h8421;
defparam \Equal2~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N23
dffeas \addr[27] (
	.clk(CLK),
	.d(\ramif.ramaddr [27]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[27]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[27] .is_wysiwyg = "true";
defparam \addr[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N17
dffeas \addr[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr22),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[26]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[26] .is_wysiwyg = "true";
defparam \addr[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N16
cycloneive_lcell_comb \Equal2~16 (
// Equation(s):
// \Equal2~16_combout  = (\ramaddr~53_combout  & (addr[27] & (addr[26] $ (!\ramaddr~55_combout )))) # (!\ramaddr~53_combout  & (!addr[27] & (addr[26] $ (!\ramaddr~55_combout ))))

	.dataa(\ramif.ramaddr [27]),
	.datab(addr[27]),
	.datac(addr[26]),
	.datad(ramaddr22),
	.cin(gnd),
	.combout(\Equal2~16_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~16 .lut_mask = 16'h9009;
defparam \Equal2~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N7
dffeas \addr[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr23),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[28]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[28] .is_wysiwyg = "true";
defparam \addr[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N5
dffeas \addr[29] (
	.clk(CLK),
	.d(\ramif.ramaddr [29]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[29]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[29] .is_wysiwyg = "true";
defparam \addr[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N6
cycloneive_lcell_comb \Equal2~17 (
// Equation(s):
// \Equal2~17_combout  = (\ramaddr~59_combout  & (addr[28] & (\ramaddr~57_combout  $ (!addr[29])))) # (!\ramaddr~59_combout  & (!addr[28] & (\ramaddr~57_combout  $ (!addr[29]))))

	.dataa(ramaddr23),
	.datab(\ramif.ramaddr [29]),
	.datac(addr[28]),
	.datad(addr[29]),
	.cin(gnd),
	.combout(\Equal2~17_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~17 .lut_mask = 16'h8421;
defparam \Equal2~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N6
cycloneive_lcell_comb \Equal2~19 (
// Equation(s):
// \Equal2~19_combout  = (\Equal2~15_combout  & (\Equal2~18_combout  & (\Equal2~16_combout  & \Equal2~17_combout )))

	.dataa(\Equal2~15_combout ),
	.datab(\Equal2~18_combout ),
	.datac(\Equal2~16_combout ),
	.datad(\Equal2~17_combout ),
	.cin(gnd),
	.combout(\Equal2~19_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~19 .lut_mask = 16'h8000;
defparam \Equal2~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N13
dffeas \addr[19] (
	.clk(CLK),
	.d(\ramif.ramaddr [19]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[19]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[19] .is_wysiwyg = "true";
defparam \addr[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y34_N11
dffeas \addr[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr17),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[18]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[18] .is_wysiwyg = "true";
defparam \addr[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N10
cycloneive_lcell_comb \Equal2~11 (
// Equation(s):
// \Equal2~11_combout  = (\ramaddr~39_combout  & (addr[18] & (addr[19] $ (!\ramaddr~37_combout )))) # (!\ramaddr~39_combout  & (!addr[18] & (addr[19] $ (!\ramaddr~37_combout ))))

	.dataa(ramaddr17),
	.datab(addr[19]),
	.datac(addr[18]),
	.datad(\ramif.ramaddr [19]),
	.cin(gnd),
	.combout(\Equal2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~11 .lut_mask = 16'h8421;
defparam \Equal2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N21
dffeas \addr[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr19),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[22]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[22] .is_wysiwyg = "true";
defparam \addr[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N20
cycloneive_lcell_comb \Equal2~13 (
// Equation(s):
// \Equal2~13_combout  = (addr[23] & (\ramaddr~45_combout  & (\ramaddr~47_combout  $ (!addr[22])))) # (!addr[23] & (!\ramaddr~45_combout  & (\ramaddr~47_combout  $ (!addr[22]))))

	.dataa(addr[23]),
	.datab(ramaddr19),
	.datac(addr[22]),
	.datad(\ramif.ramaddr [23]),
	.cin(gnd),
	.combout(\Equal2~13_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~13 .lut_mask = 16'h8241;
defparam \Equal2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N15
dffeas \addr[21] (
	.clk(CLK),
	.d(\ramif.ramaddr [21]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[21]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[21] .is_wysiwyg = "true";
defparam \addr[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N25
dffeas \addr[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr18),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[20]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[20] .is_wysiwyg = "true";
defparam \addr[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N24
cycloneive_lcell_comb \Equal2~12 (
// Equation(s):
// \Equal2~12_combout  = (\ramaddr~43_combout  & (addr[20] & (addr[21] $ (!\ramaddr~41_combout )))) # (!\ramaddr~43_combout  & (!addr[20] & (addr[21] $ (!\ramaddr~41_combout ))))

	.dataa(ramaddr18),
	.datab(addr[21]),
	.datac(addr[20]),
	.datad(\ramif.ramaddr [21]),
	.cin(gnd),
	.combout(\Equal2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~12 .lut_mask = 16'h8421;
defparam \Equal2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N18
cycloneive_lcell_comb \Equal2~14 (
// Equation(s):
// \Equal2~14_combout  = (\Equal2~10_combout  & (\Equal2~11_combout  & (\Equal2~13_combout  & \Equal2~12_combout )))

	.dataa(\Equal2~10_combout ),
	.datab(\Equal2~11_combout ),
	.datac(\Equal2~13_combout ),
	.datad(\Equal2~12_combout ),
	.cin(gnd),
	.combout(\Equal2~14_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~14 .lut_mask = 16'h8000;
defparam \Equal2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y32_N5
dffeas \addr[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr11),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[10]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[10] .is_wysiwyg = "true";
defparam \addr[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N4
cycloneive_lcell_comb \Equal2~6 (
// Equation(s):
// \Equal2~6_combout  = (addr[11] & (\ramaddr~21_combout  & (\ramaddr~23_combout  $ (!addr[10])))) # (!addr[11] & (!\ramaddr~21_combout  & (\ramaddr~23_combout  $ (!addr[10]))))

	.dataa(addr[11]),
	.datab(ramaddr11),
	.datac(addr[10]),
	.datad(ramaddr10),
	.cin(gnd),
	.combout(\Equal2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~6 .lut_mask = 16'h8241;
defparam \Equal2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y32_N1
dffeas \addr[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr9),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[8]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[8] .is_wysiwyg = "true";
defparam \addr[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N0
cycloneive_lcell_comb \Equal2~5 (
// Equation(s):
// \Equal2~5_combout  = (addr[9] & (\ramaddr~17_combout  & (addr[8] $ (!\ramaddr~19_combout )))) # (!addr[9] & (!\ramaddr~17_combout  & (addr[8] $ (!\ramaddr~19_combout ))))

	.dataa(addr[9]),
	.datab(ramaddr8),
	.datac(addr[8]),
	.datad(ramaddr9),
	.cin(gnd),
	.combout(\Equal2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~5 .lut_mask = 16'h9009;
defparam \Equal2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N25
dffeas \addr[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr15),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[14]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[14] .is_wysiwyg = "true";
defparam \addr[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N24
cycloneive_lcell_comb \Equal2~8 (
// Equation(s):
// \Equal2~8_combout  = (addr[15] & (!\ramaddr~29_combout  & (addr[14] $ (!\ramaddr~31_combout )))) # (!addr[15] & (\ramaddr~29_combout  & (addr[14] $ (!\ramaddr~31_combout ))))

	.dataa(addr[15]),
	.datab(ramaddr14),
	.datac(addr[14]),
	.datad(ramaddr15),
	.cin(gnd),
	.combout(\Equal2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~8 .lut_mask = 16'h6006;
defparam \Equal2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N8
cycloneive_lcell_comb \Equal2~9 (
// Equation(s):
// \Equal2~9_combout  = (\Equal2~7_combout  & (\Equal2~6_combout  & (\Equal2~5_combout  & \Equal2~8_combout )))

	.dataa(\Equal2~7_combout ),
	.datab(\Equal2~6_combout ),
	.datac(\Equal2~5_combout ),
	.datad(\Equal2~8_combout ),
	.cin(gnd),
	.combout(\Equal2~9_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~9 .lut_mask = 16'h8000;
defparam \Equal2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N29
dffeas \addr[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr5),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[4]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[4] .is_wysiwyg = "true";
defparam \addr[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N28
cycloneive_lcell_comb \Equal2~2 (
// Equation(s):
// \Equal2~2_combout  = (addr[5] & (\ramaddr~9_combout  & (\ramaddr~11_combout  $ (!addr[4])))) # (!addr[5] & (!\ramaddr~9_combout  & (\ramaddr~11_combout  $ (!addr[4]))))

	.dataa(addr[5]),
	.datab(ramaddr5),
	.datac(addr[4]),
	.datad(ramaddr4),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~2 .lut_mask = 16'h8241;
defparam \Equal2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y33_N3
dffeas \addr[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[1]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[1] .is_wysiwyg = "true";
defparam \addr[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N5
dffeas \addr[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr1),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[0]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[0] .is_wysiwyg = "true";
defparam \addr[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N4
cycloneive_lcell_comb \Equal2~0 (
// Equation(s):
// \Equal2~0_combout  = (\ramaddr~3_combout  & (addr[0] & (addr[1] $ (!\ramaddr~1_combout )))) # (!\ramaddr~3_combout  & (!addr[0] & (addr[1] $ (!\ramaddr~1_combout ))))

	.dataa(ramaddr1),
	.datab(addr[1]),
	.datac(addr[0]),
	.datad(ramaddr),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~0 .lut_mask = 16'h8421;
defparam \Equal2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N29
dffeas \addr[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr7),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[6]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[6] .is_wysiwyg = "true";
defparam \addr[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N28
cycloneive_lcell_comb \Equal2~3 (
// Equation(s):
// \Equal2~3_combout  = (addr[7] & (\ramaddr~13_combout  & (\ramaddr~15_combout  $ (!addr[6])))) # (!addr[7] & (!\ramaddr~13_combout  & (\ramaddr~15_combout  $ (!addr[6]))))

	.dataa(addr[7]),
	.datab(ramaddr7),
	.datac(addr[6]),
	.datad(ramaddr6),
	.cin(gnd),
	.combout(\Equal2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~3 .lut_mask = 16'h8241;
defparam \Equal2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N10
cycloneive_lcell_comb \Equal2~4 (
// Equation(s):
// \Equal2~4_combout  = (\Equal2~1_combout  & (\Equal2~2_combout  & (\Equal2~0_combout  & \Equal2~3_combout )))

	.dataa(\Equal2~1_combout ),
	.datab(\Equal2~2_combout ),
	.datac(\Equal2~0_combout ),
	.datad(\Equal2~3_combout ),
	.cin(gnd),
	.combout(\Equal2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~4 .lut_mask = 16'h8000;
defparam \Equal2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N20
cycloneive_lcell_comb \Equal2~20 (
// Equation(s):
// \Equal2~20_combout  = (\Equal2~19_combout  & (\Equal2~14_combout  & (\Equal2~9_combout  & \Equal2~4_combout )))

	.dataa(\Equal2~19_combout ),
	.datab(\Equal2~14_combout ),
	.datac(\Equal2~9_combout ),
	.datad(\Equal2~4_combout ),
	.cin(gnd),
	.combout(\Equal2~20_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~20 .lut_mask = 16'h8000;
defparam \Equal2~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N16
cycloneive_lcell_comb \ramif.ramload[16]~16 (
// Equation(s):
// \ramif.ramload[16]~16_combout  = (\nRST~input_o  & (((\ramWEN~0_combout  & \ramREN~0_combout )) # (!\Equal2~20_combout )))

	.dataa(\ramif.ramWEN ),
	.datab(\ramif.ramREN ),
	.datac(nRST),
	.datad(\Equal2~20_combout ),
	.cin(gnd),
	.combout(\ramif.ramload[16]~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[16]~16 .lut_mask = 16'h80F0;
defparam \ramif.ramload[16]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N26
cycloneive_lcell_comb \ramif.ramload[17]~18 (
// Equation(s):
// \ramif.ramload[17]~18_combout  = (\nRST~input_o  & (((\ramWEN~0_combout  & \ramREN~0_combout )) # (!\Equal2~20_combout )))

	.dataa(\ramif.ramWEN ),
	.datab(\ramif.ramREN ),
	.datac(nRST),
	.datad(\Equal2~20_combout ),
	.cin(gnd),
	.combout(\ramif.ramload[17]~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[17]~18 .lut_mask = 16'h80F0;
defparam \ramif.ramload[17]~18 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module altsyncram_1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



altsyncram_99f1 auto_generated(
	.ram_block3a32(ram_block3a32),
	.ram_block3a0(ram_block3a0),
	.ram_block3a33(ram_block3a33),
	.ram_block3a1(ram_block3a1),
	.ram_block3a34(ram_block3a34),
	.ram_block3a2(ram_block3a2),
	.ram_block3a35(ram_block3a35),
	.ram_block3a3(ram_block3a3),
	.ram_block3a36(ram_block3a36),
	.ram_block3a4(ram_block3a4),
	.ram_block3a37(ram_block3a37),
	.ram_block3a5(ram_block3a5),
	.ram_block3a38(ram_block3a38),
	.ram_block3a6(ram_block3a6),
	.ram_block3a39(ram_block3a39),
	.ram_block3a7(ram_block3a7),
	.ram_block3a40(ram_block3a40),
	.ram_block3a8(ram_block3a8),
	.ram_block3a41(ram_block3a41),
	.ram_block3a9(ram_block3a9),
	.ram_block3a42(ram_block3a42),
	.ram_block3a10(ram_block3a10),
	.ram_block3a43(ram_block3a43),
	.ram_block3a11(ram_block3a11),
	.ram_block3a44(ram_block3a44),
	.ram_block3a12(ram_block3a12),
	.ram_block3a45(ram_block3a45),
	.ram_block3a13(ram_block3a13),
	.ram_block3a46(ram_block3a46),
	.ram_block3a14(ram_block3a14),
	.ram_block3a47(ram_block3a47),
	.ram_block3a15(ram_block3a15),
	.ram_block3a48(ram_block3a48),
	.ram_block3a16(ram_block3a16),
	.ram_block3a49(ram_block3a49),
	.ram_block3a17(ram_block3a17),
	.ram_block3a50(ram_block3a50),
	.ram_block3a18(ram_block3a18),
	.ram_block3a51(ram_block3a51),
	.ram_block3a19(ram_block3a19),
	.ram_block3a52(ram_block3a52),
	.ram_block3a20(ram_block3a20),
	.ram_block3a53(ram_block3a53),
	.ram_block3a21(ram_block3a21),
	.ram_block3a54(ram_block3a54),
	.ram_block3a22(ram_block3a22),
	.ram_block3a55(ram_block3a55),
	.ram_block3a23(ram_block3a23),
	.ram_block3a56(ram_block3a56),
	.ram_block3a24(ram_block3a24),
	.ram_block3a57(ram_block3a57),
	.ram_block3a25(ram_block3a25),
	.ram_block3a58(ram_block3a58),
	.ram_block3a26(ram_block3a26),
	.ram_block3a59(ram_block3a59),
	.ram_block3a27(ram_block3a27),
	.ram_block3a60(ram_block3a60),
	.ram_block3a28(ram_block3a28),
	.ram_block3a61(ram_block3a61),
	.ram_block3a29(ram_block3a29),
	.ram_block3a62(ram_block3a62),
	.ram_block3a30(ram_block3a30),
	.ram_block3a63(ram_block3a63),
	.ram_block3a31(ram_block3a31),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.ramaddr1(ramaddr1),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_99f1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram1|ram_block3a32~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a0~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a33~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a1~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a34~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a2~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a35~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a3~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a36~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a4~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a37~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a5~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a38~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a6~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a39~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a7~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a40~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a8~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a41~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a9~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a42~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a10~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a43~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a11~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a44~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a12~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a45~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a13~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a46~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a14~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a47~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a15~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a48~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a16~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a49~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a17~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a50~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a18~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a51~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a19~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a52~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a20~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a53~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a21~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a54~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a22~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a55~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a23~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a56~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a24~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a57~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a25~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a58~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a26~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a59~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a27~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a60~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a28~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a61~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a29~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a62~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a30~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a63~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a31~PORTBDATAOUT0 ;
wire \mgl_prim2|sdr~0_combout ;
wire [0:0] \altsyncram1|address_reg_b ;
wire [31:0] \mgl_prim2|ram_rom_data_reg ;
wire [13:0] \mgl_prim2|ram_rom_addr_reg ;


sld_mod_ram_rom mgl_prim2(
	.ram_block3a32(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a0(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a33(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a1(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a34(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a2(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a35(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a3(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a36(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a4(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a37(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a5(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a38(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a6(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a39(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a7(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a40(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a8(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a41(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a9(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a42(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a10(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a43(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a11(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a44(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a12(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a45(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a13(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a46(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a14(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a47(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a15(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a48(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a16(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a49(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a17(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a50(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a18(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a51(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a19(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a52(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a20(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a53(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a21(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a54(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a22(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a55(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a23(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a56(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a24(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a57(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a25(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a58(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a26(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a59(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a27(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a60(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a28(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a61(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a29(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a62(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a30(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a63(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a31(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.is_in_use_reg1(is_in_use_reg),
	.ram_rom_data_reg_0(\mgl_prim2|ram_rom_data_reg [0]),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.ram_rom_addr_reg_0(\mgl_prim2|ram_rom_addr_reg [0]),
	.ram_rom_addr_reg_1(\mgl_prim2|ram_rom_addr_reg [1]),
	.ram_rom_addr_reg_2(\mgl_prim2|ram_rom_addr_reg [2]),
	.ram_rom_addr_reg_3(\mgl_prim2|ram_rom_addr_reg [3]),
	.ram_rom_addr_reg_4(\mgl_prim2|ram_rom_addr_reg [4]),
	.ram_rom_addr_reg_5(\mgl_prim2|ram_rom_addr_reg [5]),
	.ram_rom_addr_reg_6(\mgl_prim2|ram_rom_addr_reg [6]),
	.ram_rom_addr_reg_7(\mgl_prim2|ram_rom_addr_reg [7]),
	.ram_rom_addr_reg_8(\mgl_prim2|ram_rom_addr_reg [8]),
	.ram_rom_addr_reg_9(\mgl_prim2|ram_rom_addr_reg [9]),
	.ram_rom_addr_reg_10(\mgl_prim2|ram_rom_addr_reg [10]),
	.ram_rom_addr_reg_11(\mgl_prim2|ram_rom_addr_reg [11]),
	.ram_rom_addr_reg_12(\mgl_prim2|ram_rom_addr_reg [12]),
	.ram_rom_data_reg_1(\mgl_prim2|ram_rom_data_reg [1]),
	.ram_rom_data_reg_2(\mgl_prim2|ram_rom_data_reg [2]),
	.ram_rom_data_reg_3(\mgl_prim2|ram_rom_data_reg [3]),
	.ram_rom_data_reg_4(\mgl_prim2|ram_rom_data_reg [4]),
	.ram_rom_data_reg_5(\mgl_prim2|ram_rom_data_reg [5]),
	.ram_rom_data_reg_6(\mgl_prim2|ram_rom_data_reg [6]),
	.ram_rom_data_reg_7(\mgl_prim2|ram_rom_data_reg [7]),
	.ram_rom_data_reg_8(\mgl_prim2|ram_rom_data_reg [8]),
	.ram_rom_data_reg_9(\mgl_prim2|ram_rom_data_reg [9]),
	.ram_rom_data_reg_10(\mgl_prim2|ram_rom_data_reg [10]),
	.ram_rom_data_reg_11(\mgl_prim2|ram_rom_data_reg [11]),
	.ram_rom_data_reg_12(\mgl_prim2|ram_rom_data_reg [12]),
	.ram_rom_data_reg_13(\mgl_prim2|ram_rom_data_reg [13]),
	.ram_rom_data_reg_14(\mgl_prim2|ram_rom_data_reg [14]),
	.ram_rom_data_reg_15(\mgl_prim2|ram_rom_data_reg [15]),
	.ram_rom_data_reg_16(\mgl_prim2|ram_rom_data_reg [16]),
	.ram_rom_data_reg_17(\mgl_prim2|ram_rom_data_reg [17]),
	.ram_rom_data_reg_18(\mgl_prim2|ram_rom_data_reg [18]),
	.ram_rom_data_reg_19(\mgl_prim2|ram_rom_data_reg [19]),
	.ram_rom_data_reg_20(\mgl_prim2|ram_rom_data_reg [20]),
	.ram_rom_data_reg_21(\mgl_prim2|ram_rom_data_reg [21]),
	.ram_rom_data_reg_22(\mgl_prim2|ram_rom_data_reg [22]),
	.ram_rom_data_reg_23(\mgl_prim2|ram_rom_data_reg [23]),
	.ram_rom_data_reg_24(\mgl_prim2|ram_rom_data_reg [24]),
	.ram_rom_data_reg_25(\mgl_prim2|ram_rom_data_reg [25]),
	.ram_rom_data_reg_26(\mgl_prim2|ram_rom_data_reg [26]),
	.ram_rom_data_reg_27(\mgl_prim2|ram_rom_data_reg [27]),
	.ram_rom_data_reg_28(\mgl_prim2|ram_rom_data_reg [28]),
	.ram_rom_data_reg_29(\mgl_prim2|ram_rom_data_reg [29]),
	.ram_rom_data_reg_30(\mgl_prim2|ram_rom_data_reg [30]),
	.ram_rom_data_reg_31(\mgl_prim2|ram_rom_data_reg [31]),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.ir_in({gnd,irf_reg_3_1,gnd,gnd,irf_reg_0_1}),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.raw_tck(altera_internal_jtag1),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

altsyncram_fta2 altsyncram1(
	.ram_block3a321(ram_block3a32),
	.ram_block3a322(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a01(ram_block3a0),
	.ram_block3a02(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a331(ram_block3a33),
	.ram_block3a332(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a110(ram_block3a1),
	.ram_block3a111(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a341(ram_block3a34),
	.ram_block3a342(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a210(ram_block3a2),
	.ram_block3a211(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a351(ram_block3a35),
	.ram_block3a352(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a310(ram_block3a3),
	.ram_block3a311(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a361(ram_block3a36),
	.ram_block3a362(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a410(ram_block3a4),
	.ram_block3a411(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a371(ram_block3a37),
	.ram_block3a372(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a510(ram_block3a5),
	.ram_block3a511(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a381(ram_block3a38),
	.ram_block3a382(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a64(ram_block3a6),
	.ram_block3a65(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a391(ram_block3a39),
	.ram_block3a392(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a71(ram_block3a7),
	.ram_block3a72(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a401(ram_block3a40),
	.ram_block3a402(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a81(ram_block3a8),
	.ram_block3a82(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a412(ram_block3a41),
	.ram_block3a413(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a91(ram_block3a9),
	.ram_block3a92(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a421(ram_block3a42),
	.ram_block3a422(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a101(ram_block3a10),
	.ram_block3a102(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a431(ram_block3a43),
	.ram_block3a432(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a112(ram_block3a11),
	.ram_block3a113(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a441(ram_block3a44),
	.ram_block3a442(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a121(ram_block3a12),
	.ram_block3a122(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a451(ram_block3a45),
	.ram_block3a452(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a131(ram_block3a13),
	.ram_block3a132(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a461(ram_block3a46),
	.ram_block3a462(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a141(ram_block3a14),
	.ram_block3a142(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a471(ram_block3a47),
	.ram_block3a472(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a151(ram_block3a15),
	.ram_block3a152(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a481(ram_block3a48),
	.ram_block3a482(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a161(ram_block3a16),
	.ram_block3a162(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a491(ram_block3a49),
	.ram_block3a492(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a171(ram_block3a17),
	.ram_block3a172(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a501(ram_block3a50),
	.ram_block3a502(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a181(ram_block3a18),
	.ram_block3a182(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a512(ram_block3a51),
	.ram_block3a513(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a191(ram_block3a19),
	.ram_block3a192(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a521(ram_block3a52),
	.ram_block3a522(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a201(ram_block3a20),
	.ram_block3a202(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a531(ram_block3a53),
	.ram_block3a532(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a212(ram_block3a21),
	.ram_block3a213(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a541(ram_block3a54),
	.ram_block3a542(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a221(ram_block3a22),
	.ram_block3a222(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a551(ram_block3a55),
	.ram_block3a552(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a231(ram_block3a23),
	.ram_block3a232(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a561(ram_block3a56),
	.ram_block3a562(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a241(ram_block3a24),
	.ram_block3a242(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a571(ram_block3a57),
	.ram_block3a572(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a251(ram_block3a25),
	.ram_block3a252(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a581(ram_block3a58),
	.ram_block3a582(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a261(ram_block3a26),
	.ram_block3a262(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a591(ram_block3a59),
	.ram_block3a592(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a271(ram_block3a27),
	.ram_block3a272(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a601(ram_block3a60),
	.ram_block3a602(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a281(ram_block3a28),
	.ram_block3a282(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a611(ram_block3a61),
	.ram_block3a612(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a291(ram_block3a29),
	.ram_block3a292(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a621(ram_block3a62),
	.ram_block3a622(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a301(ram_block3a30),
	.ram_block3a302(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a631(ram_block3a63),
	.ram_block3a632(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a312(ram_block3a31),
	.ram_block3a313(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.data_b({\mgl_prim2|ram_rom_data_reg [31],\mgl_prim2|ram_rom_data_reg [30],\mgl_prim2|ram_rom_data_reg [29],\mgl_prim2|ram_rom_data_reg [28],\mgl_prim2|ram_rom_data_reg [27],\mgl_prim2|ram_rom_data_reg [26],\mgl_prim2|ram_rom_data_reg [25],\mgl_prim2|ram_rom_data_reg [24],\mgl_prim2|ram_rom_data_reg [23],
\mgl_prim2|ram_rom_data_reg [22],\mgl_prim2|ram_rom_data_reg [21],\mgl_prim2|ram_rom_data_reg [20],\mgl_prim2|ram_rom_data_reg [19],\mgl_prim2|ram_rom_data_reg [18],\mgl_prim2|ram_rom_data_reg [17],\mgl_prim2|ram_rom_data_reg [16],\mgl_prim2|ram_rom_data_reg [15],\mgl_prim2|ram_rom_data_reg [14],
\mgl_prim2|ram_rom_data_reg [13],\mgl_prim2|ram_rom_data_reg [12],\mgl_prim2|ram_rom_data_reg [11],\mgl_prim2|ram_rom_data_reg [10],\mgl_prim2|ram_rom_data_reg [9],\mgl_prim2|ram_rom_data_reg [8],\mgl_prim2|ram_rom_data_reg [7],\mgl_prim2|ram_rom_data_reg [6],\mgl_prim2|ram_rom_data_reg [5],
\mgl_prim2|ram_rom_data_reg [4],\mgl_prim2|ram_rom_data_reg [3],\mgl_prim2|ram_rom_data_reg [2],\mgl_prim2|ram_rom_data_reg [1],\mgl_prim2|ram_rom_data_reg [0]}),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.address_b({gnd,\mgl_prim2|ram_rom_addr_reg [12],\mgl_prim2|ram_rom_addr_reg [11],\mgl_prim2|ram_rom_addr_reg [10],\mgl_prim2|ram_rom_addr_reg [9],\mgl_prim2|ram_rom_addr_reg [8],\mgl_prim2|ram_rom_addr_reg [7],\mgl_prim2|ram_rom_addr_reg [6],\mgl_prim2|ram_rom_addr_reg [5],\mgl_prim2|ram_rom_addr_reg [4],
\mgl_prim2|ram_rom_addr_reg [3],\mgl_prim2|ram_rom_addr_reg [2],\mgl_prim2|ram_rom_addr_reg [1],\mgl_prim2|ram_rom_addr_reg [0]}),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.ramaddr1(ramaddr1),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.clock1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_fta2 (
	ram_block3a321,
	ram_block3a322,
	ram_block3a01,
	ram_block3a02,
	ram_block3a331,
	ram_block3a332,
	ram_block3a110,
	ram_block3a111,
	ram_block3a341,
	ram_block3a342,
	ram_block3a210,
	ram_block3a211,
	ram_block3a351,
	ram_block3a352,
	ram_block3a310,
	ram_block3a311,
	ram_block3a361,
	ram_block3a362,
	ram_block3a410,
	ram_block3a411,
	ram_block3a371,
	ram_block3a372,
	ram_block3a510,
	ram_block3a511,
	ram_block3a381,
	ram_block3a382,
	ram_block3a64,
	ram_block3a65,
	ram_block3a391,
	ram_block3a392,
	ram_block3a71,
	ram_block3a72,
	ram_block3a401,
	ram_block3a402,
	ram_block3a81,
	ram_block3a82,
	ram_block3a412,
	ram_block3a413,
	ram_block3a91,
	ram_block3a92,
	ram_block3a421,
	ram_block3a422,
	ram_block3a101,
	ram_block3a102,
	ram_block3a431,
	ram_block3a432,
	ram_block3a112,
	ram_block3a113,
	ram_block3a441,
	ram_block3a442,
	ram_block3a121,
	ram_block3a122,
	ram_block3a451,
	ram_block3a452,
	ram_block3a131,
	ram_block3a132,
	ram_block3a461,
	ram_block3a462,
	ram_block3a141,
	ram_block3a142,
	ram_block3a471,
	ram_block3a472,
	ram_block3a151,
	ram_block3a152,
	ram_block3a481,
	ram_block3a482,
	ram_block3a161,
	ram_block3a162,
	ram_block3a491,
	ram_block3a492,
	ram_block3a171,
	ram_block3a172,
	ram_block3a501,
	ram_block3a502,
	ram_block3a181,
	ram_block3a182,
	ram_block3a512,
	ram_block3a513,
	ram_block3a191,
	ram_block3a192,
	ram_block3a521,
	ram_block3a522,
	ram_block3a201,
	ram_block3a202,
	ram_block3a531,
	ram_block3a532,
	ram_block3a212,
	ram_block3a213,
	ram_block3a541,
	ram_block3a542,
	ram_block3a221,
	ram_block3a222,
	ram_block3a551,
	ram_block3a552,
	ram_block3a231,
	ram_block3a232,
	ram_block3a561,
	ram_block3a562,
	ram_block3a241,
	ram_block3a242,
	ram_block3a571,
	ram_block3a572,
	ram_block3a251,
	ram_block3a252,
	ram_block3a581,
	ram_block3a582,
	ram_block3a261,
	ram_block3a262,
	ram_block3a591,
	ram_block3a592,
	ram_block3a271,
	ram_block3a272,
	ram_block3a601,
	ram_block3a602,
	ram_block3a281,
	ram_block3a282,
	ram_block3a611,
	ram_block3a612,
	ram_block3a291,
	ram_block3a292,
	ram_block3a621,
	ram_block3a622,
	ram_block3a301,
	ram_block3a302,
	ram_block3a631,
	ram_block3a632,
	ram_block3a312,
	ram_block3a313,
	data_b,
	ram_rom_addr_reg_13,
	address_b,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	sdr,
	data_a,
	address_reg_b_0,
	ramaddr1,
	irf_reg_2_1,
	state_5,
	clock1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a321;
output 	ram_block3a322;
output 	ram_block3a01;
output 	ram_block3a02;
output 	ram_block3a331;
output 	ram_block3a332;
output 	ram_block3a110;
output 	ram_block3a111;
output 	ram_block3a341;
output 	ram_block3a342;
output 	ram_block3a210;
output 	ram_block3a211;
output 	ram_block3a351;
output 	ram_block3a352;
output 	ram_block3a310;
output 	ram_block3a311;
output 	ram_block3a361;
output 	ram_block3a362;
output 	ram_block3a410;
output 	ram_block3a411;
output 	ram_block3a371;
output 	ram_block3a372;
output 	ram_block3a510;
output 	ram_block3a511;
output 	ram_block3a381;
output 	ram_block3a382;
output 	ram_block3a64;
output 	ram_block3a65;
output 	ram_block3a391;
output 	ram_block3a392;
output 	ram_block3a71;
output 	ram_block3a72;
output 	ram_block3a401;
output 	ram_block3a402;
output 	ram_block3a81;
output 	ram_block3a82;
output 	ram_block3a412;
output 	ram_block3a413;
output 	ram_block3a91;
output 	ram_block3a92;
output 	ram_block3a421;
output 	ram_block3a422;
output 	ram_block3a101;
output 	ram_block3a102;
output 	ram_block3a431;
output 	ram_block3a432;
output 	ram_block3a112;
output 	ram_block3a113;
output 	ram_block3a441;
output 	ram_block3a442;
output 	ram_block3a121;
output 	ram_block3a122;
output 	ram_block3a451;
output 	ram_block3a452;
output 	ram_block3a131;
output 	ram_block3a132;
output 	ram_block3a461;
output 	ram_block3a462;
output 	ram_block3a141;
output 	ram_block3a142;
output 	ram_block3a471;
output 	ram_block3a472;
output 	ram_block3a151;
output 	ram_block3a152;
output 	ram_block3a481;
output 	ram_block3a482;
output 	ram_block3a161;
output 	ram_block3a162;
output 	ram_block3a491;
output 	ram_block3a492;
output 	ram_block3a171;
output 	ram_block3a172;
output 	ram_block3a501;
output 	ram_block3a502;
output 	ram_block3a181;
output 	ram_block3a182;
output 	ram_block3a512;
output 	ram_block3a513;
output 	ram_block3a191;
output 	ram_block3a192;
output 	ram_block3a521;
output 	ram_block3a522;
output 	ram_block3a201;
output 	ram_block3a202;
output 	ram_block3a531;
output 	ram_block3a532;
output 	ram_block3a212;
output 	ram_block3a213;
output 	ram_block3a541;
output 	ram_block3a542;
output 	ram_block3a221;
output 	ram_block3a222;
output 	ram_block3a551;
output 	ram_block3a552;
output 	ram_block3a231;
output 	ram_block3a232;
output 	ram_block3a561;
output 	ram_block3a562;
output 	ram_block3a241;
output 	ram_block3a242;
output 	ram_block3a571;
output 	ram_block3a572;
output 	ram_block3a251;
output 	ram_block3a252;
output 	ram_block3a581;
output 	ram_block3a582;
output 	ram_block3a261;
output 	ram_block3a262;
output 	ram_block3a591;
output 	ram_block3a592;
output 	ram_block3a271;
output 	ram_block3a272;
output 	ram_block3a601;
output 	ram_block3a602;
output 	ram_block3a281;
output 	ram_block3a282;
output 	ram_block3a611;
output 	ram_block3a612;
output 	ram_block3a291;
output 	ram_block3a292;
output 	ram_block3a621;
output 	ram_block3a622;
output 	ram_block3a301;
output 	ram_block3a302;
output 	ram_block3a631;
output 	ram_block3a632;
output 	ram_block3a312;
output 	ram_block3a313;
input 	[31:0] data_b;
input 	ram_rom_addr_reg_13;
input 	[13:0] address_b;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
input 	sdr;
input 	[31:0] data_a;
output 	address_reg_b_0;
input 	ramaddr1;
input 	irf_reg_2_1;
input 	state_5;
input 	clock1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \decode4|eq_node[1]~0_combout ;
wire \decode5|eq_node[1]~0_combout ;
wire \decode4|eq_node[0]~1_combout ;
wire \decode5|eq_node[0]~1_combout ;
wire \address_reg_b[0]~feeder_combout ;

wire [0:0] ram_block3a32_PORTADATAOUT_bus;
wire [0:0] ram_block3a32_PORTBDATAOUT_bus;
wire [0:0] ram_block3a0_PORTADATAOUT_bus;
wire [0:0] ram_block3a0_PORTBDATAOUT_bus;
wire [0:0] ram_block3a33_PORTADATAOUT_bus;
wire [0:0] ram_block3a33_PORTBDATAOUT_bus;
wire [0:0] ram_block3a1_PORTADATAOUT_bus;
wire [0:0] ram_block3a1_PORTBDATAOUT_bus;
wire [0:0] ram_block3a34_PORTADATAOUT_bus;
wire [0:0] ram_block3a34_PORTBDATAOUT_bus;
wire [0:0] ram_block3a2_PORTADATAOUT_bus;
wire [0:0] ram_block3a2_PORTBDATAOUT_bus;
wire [0:0] ram_block3a35_PORTADATAOUT_bus;
wire [0:0] ram_block3a35_PORTBDATAOUT_bus;
wire [0:0] ram_block3a3_PORTADATAOUT_bus;
wire [0:0] ram_block3a3_PORTBDATAOUT_bus;
wire [0:0] ram_block3a36_PORTADATAOUT_bus;
wire [0:0] ram_block3a36_PORTBDATAOUT_bus;
wire [0:0] ram_block3a4_PORTADATAOUT_bus;
wire [0:0] ram_block3a4_PORTBDATAOUT_bus;
wire [0:0] ram_block3a37_PORTADATAOUT_bus;
wire [0:0] ram_block3a37_PORTBDATAOUT_bus;
wire [0:0] ram_block3a5_PORTADATAOUT_bus;
wire [0:0] ram_block3a5_PORTBDATAOUT_bus;
wire [0:0] ram_block3a38_PORTADATAOUT_bus;
wire [0:0] ram_block3a38_PORTBDATAOUT_bus;
wire [0:0] ram_block3a6_PORTADATAOUT_bus;
wire [0:0] ram_block3a6_PORTBDATAOUT_bus;
wire [0:0] ram_block3a39_PORTADATAOUT_bus;
wire [0:0] ram_block3a39_PORTBDATAOUT_bus;
wire [0:0] ram_block3a7_PORTADATAOUT_bus;
wire [0:0] ram_block3a7_PORTBDATAOUT_bus;
wire [0:0] ram_block3a40_PORTADATAOUT_bus;
wire [0:0] ram_block3a40_PORTBDATAOUT_bus;
wire [0:0] ram_block3a8_PORTADATAOUT_bus;
wire [0:0] ram_block3a8_PORTBDATAOUT_bus;
wire [0:0] ram_block3a41_PORTADATAOUT_bus;
wire [0:0] ram_block3a41_PORTBDATAOUT_bus;
wire [0:0] ram_block3a9_PORTADATAOUT_bus;
wire [0:0] ram_block3a9_PORTBDATAOUT_bus;
wire [0:0] ram_block3a42_PORTADATAOUT_bus;
wire [0:0] ram_block3a42_PORTBDATAOUT_bus;
wire [0:0] ram_block3a10_PORTADATAOUT_bus;
wire [0:0] ram_block3a10_PORTBDATAOUT_bus;
wire [0:0] ram_block3a43_PORTADATAOUT_bus;
wire [0:0] ram_block3a43_PORTBDATAOUT_bus;
wire [0:0] ram_block3a11_PORTADATAOUT_bus;
wire [0:0] ram_block3a11_PORTBDATAOUT_bus;
wire [0:0] ram_block3a44_PORTADATAOUT_bus;
wire [0:0] ram_block3a44_PORTBDATAOUT_bus;
wire [0:0] ram_block3a12_PORTADATAOUT_bus;
wire [0:0] ram_block3a12_PORTBDATAOUT_bus;
wire [0:0] ram_block3a45_PORTADATAOUT_bus;
wire [0:0] ram_block3a45_PORTBDATAOUT_bus;
wire [0:0] ram_block3a13_PORTADATAOUT_bus;
wire [0:0] ram_block3a13_PORTBDATAOUT_bus;
wire [0:0] ram_block3a46_PORTADATAOUT_bus;
wire [0:0] ram_block3a46_PORTBDATAOUT_bus;
wire [0:0] ram_block3a14_PORTADATAOUT_bus;
wire [0:0] ram_block3a14_PORTBDATAOUT_bus;
wire [0:0] ram_block3a47_PORTADATAOUT_bus;
wire [0:0] ram_block3a47_PORTBDATAOUT_bus;
wire [0:0] ram_block3a15_PORTADATAOUT_bus;
wire [0:0] ram_block3a15_PORTBDATAOUT_bus;
wire [0:0] ram_block3a48_PORTADATAOUT_bus;
wire [0:0] ram_block3a48_PORTBDATAOUT_bus;
wire [0:0] ram_block3a16_PORTADATAOUT_bus;
wire [0:0] ram_block3a16_PORTBDATAOUT_bus;
wire [0:0] ram_block3a49_PORTADATAOUT_bus;
wire [0:0] ram_block3a49_PORTBDATAOUT_bus;
wire [0:0] ram_block3a17_PORTADATAOUT_bus;
wire [0:0] ram_block3a17_PORTBDATAOUT_bus;
wire [0:0] ram_block3a50_PORTADATAOUT_bus;
wire [0:0] ram_block3a50_PORTBDATAOUT_bus;
wire [0:0] ram_block3a18_PORTADATAOUT_bus;
wire [0:0] ram_block3a18_PORTBDATAOUT_bus;
wire [0:0] ram_block3a51_PORTADATAOUT_bus;
wire [0:0] ram_block3a51_PORTBDATAOUT_bus;
wire [0:0] ram_block3a19_PORTADATAOUT_bus;
wire [0:0] ram_block3a19_PORTBDATAOUT_bus;
wire [0:0] ram_block3a52_PORTADATAOUT_bus;
wire [0:0] ram_block3a52_PORTBDATAOUT_bus;
wire [0:0] ram_block3a20_PORTADATAOUT_bus;
wire [0:0] ram_block3a20_PORTBDATAOUT_bus;
wire [0:0] ram_block3a53_PORTADATAOUT_bus;
wire [0:0] ram_block3a53_PORTBDATAOUT_bus;
wire [0:0] ram_block3a21_PORTADATAOUT_bus;
wire [0:0] ram_block3a21_PORTBDATAOUT_bus;
wire [0:0] ram_block3a54_PORTADATAOUT_bus;
wire [0:0] ram_block3a54_PORTBDATAOUT_bus;
wire [0:0] ram_block3a22_PORTADATAOUT_bus;
wire [0:0] ram_block3a22_PORTBDATAOUT_bus;
wire [0:0] ram_block3a55_PORTADATAOUT_bus;
wire [0:0] ram_block3a55_PORTBDATAOUT_bus;
wire [0:0] ram_block3a23_PORTADATAOUT_bus;
wire [0:0] ram_block3a23_PORTBDATAOUT_bus;
wire [0:0] ram_block3a56_PORTADATAOUT_bus;
wire [0:0] ram_block3a56_PORTBDATAOUT_bus;
wire [0:0] ram_block3a24_PORTADATAOUT_bus;
wire [0:0] ram_block3a24_PORTBDATAOUT_bus;
wire [0:0] ram_block3a57_PORTADATAOUT_bus;
wire [0:0] ram_block3a57_PORTBDATAOUT_bus;
wire [0:0] ram_block3a25_PORTADATAOUT_bus;
wire [0:0] ram_block3a25_PORTBDATAOUT_bus;
wire [0:0] ram_block3a58_PORTADATAOUT_bus;
wire [0:0] ram_block3a58_PORTBDATAOUT_bus;
wire [0:0] ram_block3a26_PORTADATAOUT_bus;
wire [0:0] ram_block3a26_PORTBDATAOUT_bus;
wire [0:0] ram_block3a59_PORTADATAOUT_bus;
wire [0:0] ram_block3a59_PORTBDATAOUT_bus;
wire [0:0] ram_block3a27_PORTADATAOUT_bus;
wire [0:0] ram_block3a27_PORTBDATAOUT_bus;
wire [0:0] ram_block3a60_PORTADATAOUT_bus;
wire [0:0] ram_block3a60_PORTBDATAOUT_bus;
wire [0:0] ram_block3a28_PORTADATAOUT_bus;
wire [0:0] ram_block3a28_PORTBDATAOUT_bus;
wire [0:0] ram_block3a61_PORTADATAOUT_bus;
wire [0:0] ram_block3a61_PORTBDATAOUT_bus;
wire [0:0] ram_block3a29_PORTADATAOUT_bus;
wire [0:0] ram_block3a29_PORTBDATAOUT_bus;
wire [0:0] ram_block3a62_PORTADATAOUT_bus;
wire [0:0] ram_block3a62_PORTBDATAOUT_bus;
wire [0:0] ram_block3a30_PORTADATAOUT_bus;
wire [0:0] ram_block3a30_PORTBDATAOUT_bus;
wire [0:0] ram_block3a63_PORTADATAOUT_bus;
wire [0:0] ram_block3a63_PORTBDATAOUT_bus;
wire [0:0] ram_block3a31_PORTADATAOUT_bus;
wire [0:0] ram_block3a31_PORTBDATAOUT_bus;

assign ram_block3a321 = ram_block3a32_PORTADATAOUT_bus[0];

assign ram_block3a322 = ram_block3a32_PORTBDATAOUT_bus[0];

assign ram_block3a01 = ram_block3a0_PORTADATAOUT_bus[0];

assign ram_block3a02 = ram_block3a0_PORTBDATAOUT_bus[0];

assign ram_block3a331 = ram_block3a33_PORTADATAOUT_bus[0];

assign ram_block3a332 = ram_block3a33_PORTBDATAOUT_bus[0];

assign ram_block3a110 = ram_block3a1_PORTADATAOUT_bus[0];

assign ram_block3a111 = ram_block3a1_PORTBDATAOUT_bus[0];

assign ram_block3a341 = ram_block3a34_PORTADATAOUT_bus[0];

assign ram_block3a342 = ram_block3a34_PORTBDATAOUT_bus[0];

assign ram_block3a210 = ram_block3a2_PORTADATAOUT_bus[0];

assign ram_block3a211 = ram_block3a2_PORTBDATAOUT_bus[0];

assign ram_block3a351 = ram_block3a35_PORTADATAOUT_bus[0];

assign ram_block3a352 = ram_block3a35_PORTBDATAOUT_bus[0];

assign ram_block3a310 = ram_block3a3_PORTADATAOUT_bus[0];

assign ram_block3a311 = ram_block3a3_PORTBDATAOUT_bus[0];

assign ram_block3a361 = ram_block3a36_PORTADATAOUT_bus[0];

assign ram_block3a362 = ram_block3a36_PORTBDATAOUT_bus[0];

assign ram_block3a410 = ram_block3a4_PORTADATAOUT_bus[0];

assign ram_block3a411 = ram_block3a4_PORTBDATAOUT_bus[0];

assign ram_block3a371 = ram_block3a37_PORTADATAOUT_bus[0];

assign ram_block3a372 = ram_block3a37_PORTBDATAOUT_bus[0];

assign ram_block3a510 = ram_block3a5_PORTADATAOUT_bus[0];

assign ram_block3a511 = ram_block3a5_PORTBDATAOUT_bus[0];

assign ram_block3a381 = ram_block3a38_PORTADATAOUT_bus[0];

assign ram_block3a382 = ram_block3a38_PORTBDATAOUT_bus[0];

assign ram_block3a64 = ram_block3a6_PORTADATAOUT_bus[0];

assign ram_block3a65 = ram_block3a6_PORTBDATAOUT_bus[0];

assign ram_block3a391 = ram_block3a39_PORTADATAOUT_bus[0];

assign ram_block3a392 = ram_block3a39_PORTBDATAOUT_bus[0];

assign ram_block3a71 = ram_block3a7_PORTADATAOUT_bus[0];

assign ram_block3a72 = ram_block3a7_PORTBDATAOUT_bus[0];

assign ram_block3a401 = ram_block3a40_PORTADATAOUT_bus[0];

assign ram_block3a402 = ram_block3a40_PORTBDATAOUT_bus[0];

assign ram_block3a81 = ram_block3a8_PORTADATAOUT_bus[0];

assign ram_block3a82 = ram_block3a8_PORTBDATAOUT_bus[0];

assign ram_block3a412 = ram_block3a41_PORTADATAOUT_bus[0];

assign ram_block3a413 = ram_block3a41_PORTBDATAOUT_bus[0];

assign ram_block3a91 = ram_block3a9_PORTADATAOUT_bus[0];

assign ram_block3a92 = ram_block3a9_PORTBDATAOUT_bus[0];

assign ram_block3a421 = ram_block3a42_PORTADATAOUT_bus[0];

assign ram_block3a422 = ram_block3a42_PORTBDATAOUT_bus[0];

assign ram_block3a101 = ram_block3a10_PORTADATAOUT_bus[0];

assign ram_block3a102 = ram_block3a10_PORTBDATAOUT_bus[0];

assign ram_block3a431 = ram_block3a43_PORTADATAOUT_bus[0];

assign ram_block3a432 = ram_block3a43_PORTBDATAOUT_bus[0];

assign ram_block3a112 = ram_block3a11_PORTADATAOUT_bus[0];

assign ram_block3a113 = ram_block3a11_PORTBDATAOUT_bus[0];

assign ram_block3a441 = ram_block3a44_PORTADATAOUT_bus[0];

assign ram_block3a442 = ram_block3a44_PORTBDATAOUT_bus[0];

assign ram_block3a121 = ram_block3a12_PORTADATAOUT_bus[0];

assign ram_block3a122 = ram_block3a12_PORTBDATAOUT_bus[0];

assign ram_block3a451 = ram_block3a45_PORTADATAOUT_bus[0];

assign ram_block3a452 = ram_block3a45_PORTBDATAOUT_bus[0];

assign ram_block3a131 = ram_block3a13_PORTADATAOUT_bus[0];

assign ram_block3a132 = ram_block3a13_PORTBDATAOUT_bus[0];

assign ram_block3a461 = ram_block3a46_PORTADATAOUT_bus[0];

assign ram_block3a462 = ram_block3a46_PORTBDATAOUT_bus[0];

assign ram_block3a141 = ram_block3a14_PORTADATAOUT_bus[0];

assign ram_block3a142 = ram_block3a14_PORTBDATAOUT_bus[0];

assign ram_block3a471 = ram_block3a47_PORTADATAOUT_bus[0];

assign ram_block3a472 = ram_block3a47_PORTBDATAOUT_bus[0];

assign ram_block3a151 = ram_block3a15_PORTADATAOUT_bus[0];

assign ram_block3a152 = ram_block3a15_PORTBDATAOUT_bus[0];

assign ram_block3a481 = ram_block3a48_PORTADATAOUT_bus[0];

assign ram_block3a482 = ram_block3a48_PORTBDATAOUT_bus[0];

assign ram_block3a161 = ram_block3a16_PORTADATAOUT_bus[0];

assign ram_block3a162 = ram_block3a16_PORTBDATAOUT_bus[0];

assign ram_block3a491 = ram_block3a49_PORTADATAOUT_bus[0];

assign ram_block3a492 = ram_block3a49_PORTBDATAOUT_bus[0];

assign ram_block3a171 = ram_block3a17_PORTADATAOUT_bus[0];

assign ram_block3a172 = ram_block3a17_PORTBDATAOUT_bus[0];

assign ram_block3a501 = ram_block3a50_PORTADATAOUT_bus[0];

assign ram_block3a502 = ram_block3a50_PORTBDATAOUT_bus[0];

assign ram_block3a181 = ram_block3a18_PORTADATAOUT_bus[0];

assign ram_block3a182 = ram_block3a18_PORTBDATAOUT_bus[0];

assign ram_block3a512 = ram_block3a51_PORTADATAOUT_bus[0];

assign ram_block3a513 = ram_block3a51_PORTBDATAOUT_bus[0];

assign ram_block3a191 = ram_block3a19_PORTADATAOUT_bus[0];

assign ram_block3a192 = ram_block3a19_PORTBDATAOUT_bus[0];

assign ram_block3a521 = ram_block3a52_PORTADATAOUT_bus[0];

assign ram_block3a522 = ram_block3a52_PORTBDATAOUT_bus[0];

assign ram_block3a201 = ram_block3a20_PORTADATAOUT_bus[0];

assign ram_block3a202 = ram_block3a20_PORTBDATAOUT_bus[0];

assign ram_block3a531 = ram_block3a53_PORTADATAOUT_bus[0];

assign ram_block3a532 = ram_block3a53_PORTBDATAOUT_bus[0];

assign ram_block3a212 = ram_block3a21_PORTADATAOUT_bus[0];

assign ram_block3a213 = ram_block3a21_PORTBDATAOUT_bus[0];

assign ram_block3a541 = ram_block3a54_PORTADATAOUT_bus[0];

assign ram_block3a542 = ram_block3a54_PORTBDATAOUT_bus[0];

assign ram_block3a221 = ram_block3a22_PORTADATAOUT_bus[0];

assign ram_block3a222 = ram_block3a22_PORTBDATAOUT_bus[0];

assign ram_block3a551 = ram_block3a55_PORTADATAOUT_bus[0];

assign ram_block3a552 = ram_block3a55_PORTBDATAOUT_bus[0];

assign ram_block3a231 = ram_block3a23_PORTADATAOUT_bus[0];

assign ram_block3a232 = ram_block3a23_PORTBDATAOUT_bus[0];

assign ram_block3a561 = ram_block3a56_PORTADATAOUT_bus[0];

assign ram_block3a562 = ram_block3a56_PORTBDATAOUT_bus[0];

assign ram_block3a241 = ram_block3a24_PORTADATAOUT_bus[0];

assign ram_block3a242 = ram_block3a24_PORTBDATAOUT_bus[0];

assign ram_block3a571 = ram_block3a57_PORTADATAOUT_bus[0];

assign ram_block3a572 = ram_block3a57_PORTBDATAOUT_bus[0];

assign ram_block3a251 = ram_block3a25_PORTADATAOUT_bus[0];

assign ram_block3a252 = ram_block3a25_PORTBDATAOUT_bus[0];

assign ram_block3a581 = ram_block3a58_PORTADATAOUT_bus[0];

assign ram_block3a582 = ram_block3a58_PORTBDATAOUT_bus[0];

assign ram_block3a261 = ram_block3a26_PORTADATAOUT_bus[0];

assign ram_block3a262 = ram_block3a26_PORTBDATAOUT_bus[0];

assign ram_block3a591 = ram_block3a59_PORTADATAOUT_bus[0];

assign ram_block3a592 = ram_block3a59_PORTBDATAOUT_bus[0];

assign ram_block3a271 = ram_block3a27_PORTADATAOUT_bus[0];

assign ram_block3a272 = ram_block3a27_PORTBDATAOUT_bus[0];

assign ram_block3a601 = ram_block3a60_PORTADATAOUT_bus[0];

assign ram_block3a602 = ram_block3a60_PORTBDATAOUT_bus[0];

assign ram_block3a281 = ram_block3a28_PORTADATAOUT_bus[0];

assign ram_block3a282 = ram_block3a28_PORTBDATAOUT_bus[0];

assign ram_block3a611 = ram_block3a61_PORTADATAOUT_bus[0];

assign ram_block3a612 = ram_block3a61_PORTBDATAOUT_bus[0];

assign ram_block3a291 = ram_block3a29_PORTADATAOUT_bus[0];

assign ram_block3a292 = ram_block3a29_PORTBDATAOUT_bus[0];

assign ram_block3a621 = ram_block3a62_PORTADATAOUT_bus[0];

assign ram_block3a622 = ram_block3a62_PORTBDATAOUT_bus[0];

assign ram_block3a301 = ram_block3a30_PORTADATAOUT_bus[0];

assign ram_block3a302 = ram_block3a30_PORTBDATAOUT_bus[0];

assign ram_block3a631 = ram_block3a63_PORTADATAOUT_bus[0];

assign ram_block3a632 = ram_block3a63_PORTBDATAOUT_bus[0];

assign ram_block3a312 = ram_block3a31_PORTADATAOUT_bus[0];

assign ram_block3a313 = ram_block3a31_PORTBDATAOUT_bus[0];

decode_jsa_1 decode5(
	.ram_rom_addr_reg_13(ram_rom_addr_reg_13),
	.sdr(sdr),
	.eq_node_1(\decode5|eq_node[1]~0_combout ),
	.eq_node_0(\decode5|eq_node[0]~1_combout ),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

decode_jsa decode4(
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.eq_node_1(\decode4|eq_node[1]~0_combout ),
	.eq_node_0(\decode4|eq_node[0]~1_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: M9K_X64_Y32_N0
cycloneive_ram_block ram_block3a32(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a32_PORTADATAOUT_bus),
	.portbdataout(ram_block3a32_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a32.clk0_core_clock_enable = "ena0";
defparam ram_block3a32.clk1_core_clock_enable = "ena1";
defparam ram_block3a32.data_interleave_offset_in_bits = 1;
defparam ram_block3a32.data_interleave_width_in_bits = 1;
defparam ram_block3a32.init_file = "meminit.hex";
defparam ram_block3a32.init_file_layout = "port_a";
defparam ram_block3a32.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a32.operation_mode = "bidir_dual_port";
defparam ram_block3a32.port_a_address_clear = "none";
defparam ram_block3a32.port_a_address_width = 13;
defparam ram_block3a32.port_a_byte_enable_clock = "none";
defparam ram_block3a32.port_a_data_out_clear = "none";
defparam ram_block3a32.port_a_data_out_clock = "none";
defparam ram_block3a32.port_a_data_width = 1;
defparam ram_block3a32.port_a_first_address = 0;
defparam ram_block3a32.port_a_first_bit_number = 0;
defparam ram_block3a32.port_a_last_address = 8191;
defparam ram_block3a32.port_a_logical_ram_depth = 16384;
defparam ram_block3a32.port_a_logical_ram_width = 32;
defparam ram_block3a32.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_address_clear = "none";
defparam ram_block3a32.port_b_address_clock = "clock1";
defparam ram_block3a32.port_b_address_width = 13;
defparam ram_block3a32.port_b_data_in_clock = "clock1";
defparam ram_block3a32.port_b_data_out_clear = "none";
defparam ram_block3a32.port_b_data_out_clock = "none";
defparam ram_block3a32.port_b_data_width = 1;
defparam ram_block3a32.port_b_first_address = 0;
defparam ram_block3a32.port_b_first_bit_number = 0;
defparam ram_block3a32.port_b_last_address = 8191;
defparam ram_block3a32.port_b_logical_ram_depth = 16384;
defparam ram_block3a32.port_b_logical_ram_width = 32;
defparam ram_block3a32.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_read_enable_clock = "clock1";
defparam ram_block3a32.port_b_write_enable_clock = "clock1";
defparam ram_block3a32.ram_block_type = "M9K";
defparam ram_block3a32.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y48_N0
cycloneive_ram_block ram_block3a0(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a0_PORTADATAOUT_bus),
	.portbdataout(ram_block3a0_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a0.clk0_core_clock_enable = "ena0";
defparam ram_block3a0.clk1_core_clock_enable = "ena1";
defparam ram_block3a0.data_interleave_offset_in_bits = 1;
defparam ram_block3a0.data_interleave_width_in_bits = 1;
defparam ram_block3a0.init_file = "meminit.hex";
defparam ram_block3a0.init_file_layout = "port_a";
defparam ram_block3a0.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a0.operation_mode = "bidir_dual_port";
defparam ram_block3a0.port_a_address_clear = "none";
defparam ram_block3a0.port_a_address_width = 13;
defparam ram_block3a0.port_a_byte_enable_clock = "none";
defparam ram_block3a0.port_a_data_out_clear = "none";
defparam ram_block3a0.port_a_data_out_clock = "none";
defparam ram_block3a0.port_a_data_width = 1;
defparam ram_block3a0.port_a_first_address = 0;
defparam ram_block3a0.port_a_first_bit_number = 0;
defparam ram_block3a0.port_a_last_address = 8191;
defparam ram_block3a0.port_a_logical_ram_depth = 16384;
defparam ram_block3a0.port_a_logical_ram_width = 32;
defparam ram_block3a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_address_clear = "none";
defparam ram_block3a0.port_b_address_clock = "clock1";
defparam ram_block3a0.port_b_address_width = 13;
defparam ram_block3a0.port_b_data_in_clock = "clock1";
defparam ram_block3a0.port_b_data_out_clear = "none";
defparam ram_block3a0.port_b_data_out_clock = "none";
defparam ram_block3a0.port_b_data_width = 1;
defparam ram_block3a0.port_b_first_address = 0;
defparam ram_block3a0.port_b_first_bit_number = 0;
defparam ram_block3a0.port_b_last_address = 8191;
defparam ram_block3a0.port_b_logical_ram_depth = 16384;
defparam ram_block3a0.port_b_logical_ram_width = 32;
defparam ram_block3a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_read_enable_clock = "clock1";
defparam ram_block3a0.port_b_write_enable_clock = "clock1";
defparam ram_block3a0.ram_block_type = "M9K";
defparam ram_block3a0.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010014AD3;
// synopsys translate_on

// Location: M9K_X64_Y49_N0
cycloneive_ram_block ram_block3a33(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a33_PORTADATAOUT_bus),
	.portbdataout(ram_block3a33_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a33.clk0_core_clock_enable = "ena0";
defparam ram_block3a33.clk1_core_clock_enable = "ena1";
defparam ram_block3a33.data_interleave_offset_in_bits = 1;
defparam ram_block3a33.data_interleave_width_in_bits = 1;
defparam ram_block3a33.init_file = "meminit.hex";
defparam ram_block3a33.init_file_layout = "port_a";
defparam ram_block3a33.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a33.operation_mode = "bidir_dual_port";
defparam ram_block3a33.port_a_address_clear = "none";
defparam ram_block3a33.port_a_address_width = 13;
defparam ram_block3a33.port_a_byte_enable_clock = "none";
defparam ram_block3a33.port_a_data_out_clear = "none";
defparam ram_block3a33.port_a_data_out_clock = "none";
defparam ram_block3a33.port_a_data_width = 1;
defparam ram_block3a33.port_a_first_address = 0;
defparam ram_block3a33.port_a_first_bit_number = 1;
defparam ram_block3a33.port_a_last_address = 8191;
defparam ram_block3a33.port_a_logical_ram_depth = 16384;
defparam ram_block3a33.port_a_logical_ram_width = 32;
defparam ram_block3a33.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_address_clear = "none";
defparam ram_block3a33.port_b_address_clock = "clock1";
defparam ram_block3a33.port_b_address_width = 13;
defparam ram_block3a33.port_b_data_in_clock = "clock1";
defparam ram_block3a33.port_b_data_out_clear = "none";
defparam ram_block3a33.port_b_data_out_clock = "none";
defparam ram_block3a33.port_b_data_width = 1;
defparam ram_block3a33.port_b_first_address = 0;
defparam ram_block3a33.port_b_first_bit_number = 1;
defparam ram_block3a33.port_b_last_address = 8191;
defparam ram_block3a33.port_b_logical_ram_depth = 16384;
defparam ram_block3a33.port_b_logical_ram_width = 32;
defparam ram_block3a33.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_read_enable_clock = "clock1";
defparam ram_block3a33.port_b_write_enable_clock = "clock1";
defparam ram_block3a33.ram_block_type = "M9K";
defparam ram_block3a33.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y34_N0
cycloneive_ram_block ram_block3a1(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a1_PORTADATAOUT_bus),
	.portbdataout(ram_block3a1_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a1.clk0_core_clock_enable = "ena0";
defparam ram_block3a1.clk1_core_clock_enable = "ena1";
defparam ram_block3a1.data_interleave_offset_in_bits = 1;
defparam ram_block3a1.data_interleave_width_in_bits = 1;
defparam ram_block3a1.init_file = "meminit.hex";
defparam ram_block3a1.init_file_layout = "port_a";
defparam ram_block3a1.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a1.operation_mode = "bidir_dual_port";
defparam ram_block3a1.port_a_address_clear = "none";
defparam ram_block3a1.port_a_address_width = 13;
defparam ram_block3a1.port_a_byte_enable_clock = "none";
defparam ram_block3a1.port_a_data_out_clear = "none";
defparam ram_block3a1.port_a_data_out_clock = "none";
defparam ram_block3a1.port_a_data_width = 1;
defparam ram_block3a1.port_a_first_address = 0;
defparam ram_block3a1.port_a_first_bit_number = 1;
defparam ram_block3a1.port_a_last_address = 8191;
defparam ram_block3a1.port_a_logical_ram_depth = 16384;
defparam ram_block3a1.port_a_logical_ram_width = 32;
defparam ram_block3a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_address_clear = "none";
defparam ram_block3a1.port_b_address_clock = "clock1";
defparam ram_block3a1.port_b_address_width = 13;
defparam ram_block3a1.port_b_data_in_clock = "clock1";
defparam ram_block3a1.port_b_data_out_clear = "none";
defparam ram_block3a1.port_b_data_out_clock = "none";
defparam ram_block3a1.port_b_data_width = 1;
defparam ram_block3a1.port_b_first_address = 0;
defparam ram_block3a1.port_b_first_bit_number = 1;
defparam ram_block3a1.port_b_last_address = 8191;
defparam ram_block3a1.port_b_logical_ram_depth = 16384;
defparam ram_block3a1.port_b_logical_ram_width = 32;
defparam ram_block3a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_read_enable_clock = "clock1";
defparam ram_block3a1.port_b_write_enable_clock = "clock1";
defparam ram_block3a1.ram_block_type = "M9K";
defparam ram_block3a1.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010018E40;
// synopsys translate_on

// Location: M9K_X37_Y32_N0
cycloneive_ram_block ram_block3a34(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a34_PORTADATAOUT_bus),
	.portbdataout(ram_block3a34_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a34.clk0_core_clock_enable = "ena0";
defparam ram_block3a34.clk1_core_clock_enable = "ena1";
defparam ram_block3a34.data_interleave_offset_in_bits = 1;
defparam ram_block3a34.data_interleave_width_in_bits = 1;
defparam ram_block3a34.init_file = "meminit.hex";
defparam ram_block3a34.init_file_layout = "port_a";
defparam ram_block3a34.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a34.operation_mode = "bidir_dual_port";
defparam ram_block3a34.port_a_address_clear = "none";
defparam ram_block3a34.port_a_address_width = 13;
defparam ram_block3a34.port_a_byte_enable_clock = "none";
defparam ram_block3a34.port_a_data_out_clear = "none";
defparam ram_block3a34.port_a_data_out_clock = "none";
defparam ram_block3a34.port_a_data_width = 1;
defparam ram_block3a34.port_a_first_address = 0;
defparam ram_block3a34.port_a_first_bit_number = 2;
defparam ram_block3a34.port_a_last_address = 8191;
defparam ram_block3a34.port_a_logical_ram_depth = 16384;
defparam ram_block3a34.port_a_logical_ram_width = 32;
defparam ram_block3a34.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_address_clear = "none";
defparam ram_block3a34.port_b_address_clock = "clock1";
defparam ram_block3a34.port_b_address_width = 13;
defparam ram_block3a34.port_b_data_in_clock = "clock1";
defparam ram_block3a34.port_b_data_out_clear = "none";
defparam ram_block3a34.port_b_data_out_clock = "none";
defparam ram_block3a34.port_b_data_width = 1;
defparam ram_block3a34.port_b_first_address = 0;
defparam ram_block3a34.port_b_first_bit_number = 2;
defparam ram_block3a34.port_b_last_address = 8191;
defparam ram_block3a34.port_b_logical_ram_depth = 16384;
defparam ram_block3a34.port_b_logical_ram_width = 32;
defparam ram_block3a34.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_read_enable_clock = "clock1";
defparam ram_block3a34.port_b_write_enable_clock = "clock1";
defparam ram_block3a34.ram_block_type = "M9K";
defparam ram_block3a34.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y29_N0
cycloneive_ram_block ram_block3a2(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a2_PORTADATAOUT_bus),
	.portbdataout(ram_block3a2_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a2.clk0_core_clock_enable = "ena0";
defparam ram_block3a2.clk1_core_clock_enable = "ena1";
defparam ram_block3a2.data_interleave_offset_in_bits = 1;
defparam ram_block3a2.data_interleave_width_in_bits = 1;
defparam ram_block3a2.init_file = "meminit.hex";
defparam ram_block3a2.init_file_layout = "port_a";
defparam ram_block3a2.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a2.operation_mode = "bidir_dual_port";
defparam ram_block3a2.port_a_address_clear = "none";
defparam ram_block3a2.port_a_address_width = 13;
defparam ram_block3a2.port_a_byte_enable_clock = "none";
defparam ram_block3a2.port_a_data_out_clear = "none";
defparam ram_block3a2.port_a_data_out_clock = "none";
defparam ram_block3a2.port_a_data_width = 1;
defparam ram_block3a2.port_a_first_address = 0;
defparam ram_block3a2.port_a_first_bit_number = 2;
defparam ram_block3a2.port_a_last_address = 8191;
defparam ram_block3a2.port_a_logical_ram_depth = 16384;
defparam ram_block3a2.port_a_logical_ram_width = 32;
defparam ram_block3a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_address_clear = "none";
defparam ram_block3a2.port_b_address_clock = "clock1";
defparam ram_block3a2.port_b_address_width = 13;
defparam ram_block3a2.port_b_data_in_clock = "clock1";
defparam ram_block3a2.port_b_data_out_clear = "none";
defparam ram_block3a2.port_b_data_out_clock = "none";
defparam ram_block3a2.port_b_data_width = 1;
defparam ram_block3a2.port_b_first_address = 0;
defparam ram_block3a2.port_b_first_bit_number = 2;
defparam ram_block3a2.port_b_last_address = 8191;
defparam ram_block3a2.port_b_logical_ram_depth = 16384;
defparam ram_block3a2.port_b_logical_ram_width = 32;
defparam ram_block3a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_read_enable_clock = "clock1";
defparam ram_block3a2.port_b_write_enable_clock = "clock1";
defparam ram_block3a2.ram_block_type = "M9K";
defparam ram_block3a2.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001AA9FC70;
// synopsys translate_on

// Location: M9K_X51_Y29_N0
cycloneive_ram_block ram_block3a35(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a35_PORTADATAOUT_bus),
	.portbdataout(ram_block3a35_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a35.clk0_core_clock_enable = "ena0";
defparam ram_block3a35.clk1_core_clock_enable = "ena1";
defparam ram_block3a35.data_interleave_offset_in_bits = 1;
defparam ram_block3a35.data_interleave_width_in_bits = 1;
defparam ram_block3a35.init_file = "meminit.hex";
defparam ram_block3a35.init_file_layout = "port_a";
defparam ram_block3a35.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a35.operation_mode = "bidir_dual_port";
defparam ram_block3a35.port_a_address_clear = "none";
defparam ram_block3a35.port_a_address_width = 13;
defparam ram_block3a35.port_a_byte_enable_clock = "none";
defparam ram_block3a35.port_a_data_out_clear = "none";
defparam ram_block3a35.port_a_data_out_clock = "none";
defparam ram_block3a35.port_a_data_width = 1;
defparam ram_block3a35.port_a_first_address = 0;
defparam ram_block3a35.port_a_first_bit_number = 3;
defparam ram_block3a35.port_a_last_address = 8191;
defparam ram_block3a35.port_a_logical_ram_depth = 16384;
defparam ram_block3a35.port_a_logical_ram_width = 32;
defparam ram_block3a35.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_address_clear = "none";
defparam ram_block3a35.port_b_address_clock = "clock1";
defparam ram_block3a35.port_b_address_width = 13;
defparam ram_block3a35.port_b_data_in_clock = "clock1";
defparam ram_block3a35.port_b_data_out_clear = "none";
defparam ram_block3a35.port_b_data_out_clock = "none";
defparam ram_block3a35.port_b_data_width = 1;
defparam ram_block3a35.port_b_first_address = 0;
defparam ram_block3a35.port_b_first_bit_number = 3;
defparam ram_block3a35.port_b_last_address = 8191;
defparam ram_block3a35.port_b_logical_ram_depth = 16384;
defparam ram_block3a35.port_b_logical_ram_width = 32;
defparam ram_block3a35.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_read_enable_clock = "clock1";
defparam ram_block3a35.port_b_write_enable_clock = "clock1";
defparam ram_block3a35.ram_block_type = "M9K";
defparam ram_block3a35.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y35_N0
cycloneive_ram_block ram_block3a3(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a3_PORTADATAOUT_bus),
	.portbdataout(ram_block3a3_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a3.clk0_core_clock_enable = "ena0";
defparam ram_block3a3.clk1_core_clock_enable = "ena1";
defparam ram_block3a3.data_interleave_offset_in_bits = 1;
defparam ram_block3a3.data_interleave_width_in_bits = 1;
defparam ram_block3a3.init_file = "meminit.hex";
defparam ram_block3a3.init_file_layout = "port_a";
defparam ram_block3a3.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a3.operation_mode = "bidir_dual_port";
defparam ram_block3a3.port_a_address_clear = "none";
defparam ram_block3a3.port_a_address_width = 13;
defparam ram_block3a3.port_a_byte_enable_clock = "none";
defparam ram_block3a3.port_a_data_out_clear = "none";
defparam ram_block3a3.port_a_data_out_clock = "none";
defparam ram_block3a3.port_a_data_width = 1;
defparam ram_block3a3.port_a_first_address = 0;
defparam ram_block3a3.port_a_first_bit_number = 3;
defparam ram_block3a3.port_a_last_address = 8191;
defparam ram_block3a3.port_a_logical_ram_depth = 16384;
defparam ram_block3a3.port_a_logical_ram_width = 32;
defparam ram_block3a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_address_clear = "none";
defparam ram_block3a3.port_b_address_clock = "clock1";
defparam ram_block3a3.port_b_address_width = 13;
defparam ram_block3a3.port_b_data_in_clock = "clock1";
defparam ram_block3a3.port_b_data_out_clear = "none";
defparam ram_block3a3.port_b_data_out_clock = "none";
defparam ram_block3a3.port_b_data_width = 1;
defparam ram_block3a3.port_b_first_address = 0;
defparam ram_block3a3.port_b_first_bit_number = 3;
defparam ram_block3a3.port_b_last_address = 8191;
defparam ram_block3a3.port_b_logical_ram_depth = 16384;
defparam ram_block3a3.port_b_logical_ram_width = 32;
defparam ram_block3a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_read_enable_clock = "clock1";
defparam ram_block3a3.port_b_write_enable_clock = "clock1";
defparam ram_block3a3.ram_block_type = "M9K";
defparam ram_block3a3.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013300841;
// synopsys translate_on

// Location: M9K_X37_Y38_N0
cycloneive_ram_block ram_block3a36(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a36_PORTADATAOUT_bus),
	.portbdataout(ram_block3a36_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a36.clk0_core_clock_enable = "ena0";
defparam ram_block3a36.clk1_core_clock_enable = "ena1";
defparam ram_block3a36.data_interleave_offset_in_bits = 1;
defparam ram_block3a36.data_interleave_width_in_bits = 1;
defparam ram_block3a36.init_file = "meminit.hex";
defparam ram_block3a36.init_file_layout = "port_a";
defparam ram_block3a36.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a36.operation_mode = "bidir_dual_port";
defparam ram_block3a36.port_a_address_clear = "none";
defparam ram_block3a36.port_a_address_width = 13;
defparam ram_block3a36.port_a_byte_enable_clock = "none";
defparam ram_block3a36.port_a_data_out_clear = "none";
defparam ram_block3a36.port_a_data_out_clock = "none";
defparam ram_block3a36.port_a_data_width = 1;
defparam ram_block3a36.port_a_first_address = 0;
defparam ram_block3a36.port_a_first_bit_number = 4;
defparam ram_block3a36.port_a_last_address = 8191;
defparam ram_block3a36.port_a_logical_ram_depth = 16384;
defparam ram_block3a36.port_a_logical_ram_width = 32;
defparam ram_block3a36.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_address_clear = "none";
defparam ram_block3a36.port_b_address_clock = "clock1";
defparam ram_block3a36.port_b_address_width = 13;
defparam ram_block3a36.port_b_data_in_clock = "clock1";
defparam ram_block3a36.port_b_data_out_clear = "none";
defparam ram_block3a36.port_b_data_out_clock = "none";
defparam ram_block3a36.port_b_data_width = 1;
defparam ram_block3a36.port_b_first_address = 0;
defparam ram_block3a36.port_b_first_bit_number = 4;
defparam ram_block3a36.port_b_last_address = 8191;
defparam ram_block3a36.port_b_logical_ram_depth = 16384;
defparam ram_block3a36.port_b_logical_ram_width = 32;
defparam ram_block3a36.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_read_enable_clock = "clock1";
defparam ram_block3a36.port_b_write_enable_clock = "clock1";
defparam ram_block3a36.ram_block_type = "M9K";
defparam ram_block3a36.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y39_N0
cycloneive_ram_block ram_block3a4(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a4_PORTADATAOUT_bus),
	.portbdataout(ram_block3a4_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a4.clk0_core_clock_enable = "ena0";
defparam ram_block3a4.clk1_core_clock_enable = "ena1";
defparam ram_block3a4.data_interleave_offset_in_bits = 1;
defparam ram_block3a4.data_interleave_width_in_bits = 1;
defparam ram_block3a4.init_file = "meminit.hex";
defparam ram_block3a4.init_file_layout = "port_a";
defparam ram_block3a4.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a4.operation_mode = "bidir_dual_port";
defparam ram_block3a4.port_a_address_clear = "none";
defparam ram_block3a4.port_a_address_width = 13;
defparam ram_block3a4.port_a_byte_enable_clock = "none";
defparam ram_block3a4.port_a_data_out_clear = "none";
defparam ram_block3a4.port_a_data_out_clock = "none";
defparam ram_block3a4.port_a_data_width = 1;
defparam ram_block3a4.port_a_first_address = 0;
defparam ram_block3a4.port_a_first_bit_number = 4;
defparam ram_block3a4.port_a_last_address = 8191;
defparam ram_block3a4.port_a_logical_ram_depth = 16384;
defparam ram_block3a4.port_a_logical_ram_width = 32;
defparam ram_block3a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_address_clear = "none";
defparam ram_block3a4.port_b_address_clock = "clock1";
defparam ram_block3a4.port_b_address_width = 13;
defparam ram_block3a4.port_b_data_in_clock = "clock1";
defparam ram_block3a4.port_b_data_out_clear = "none";
defparam ram_block3a4.port_b_data_out_clock = "none";
defparam ram_block3a4.port_b_data_width = 1;
defparam ram_block3a4.port_b_first_address = 0;
defparam ram_block3a4.port_b_first_bit_number = 4;
defparam ram_block3a4.port_b_last_address = 8191;
defparam ram_block3a4.port_b_logical_ram_depth = 16384;
defparam ram_block3a4.port_b_logical_ram_width = 32;
defparam ram_block3a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_read_enable_clock = "clock1";
defparam ram_block3a4.port_b_write_enable_clock = "clock1";
defparam ram_block3a4.ram_block_type = "M9K";
defparam ram_block3a4.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013C0080A;
// synopsys translate_on

// Location: M9K_X78_Y32_N0
cycloneive_ram_block ram_block3a37(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a37_PORTADATAOUT_bus),
	.portbdataout(ram_block3a37_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a37.clk0_core_clock_enable = "ena0";
defparam ram_block3a37.clk1_core_clock_enable = "ena1";
defparam ram_block3a37.data_interleave_offset_in_bits = 1;
defparam ram_block3a37.data_interleave_width_in_bits = 1;
defparam ram_block3a37.init_file = "meminit.hex";
defparam ram_block3a37.init_file_layout = "port_a";
defparam ram_block3a37.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a37.operation_mode = "bidir_dual_port";
defparam ram_block3a37.port_a_address_clear = "none";
defparam ram_block3a37.port_a_address_width = 13;
defparam ram_block3a37.port_a_byte_enable_clock = "none";
defparam ram_block3a37.port_a_data_out_clear = "none";
defparam ram_block3a37.port_a_data_out_clock = "none";
defparam ram_block3a37.port_a_data_width = 1;
defparam ram_block3a37.port_a_first_address = 0;
defparam ram_block3a37.port_a_first_bit_number = 5;
defparam ram_block3a37.port_a_last_address = 8191;
defparam ram_block3a37.port_a_logical_ram_depth = 16384;
defparam ram_block3a37.port_a_logical_ram_width = 32;
defparam ram_block3a37.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_address_clear = "none";
defparam ram_block3a37.port_b_address_clock = "clock1";
defparam ram_block3a37.port_b_address_width = 13;
defparam ram_block3a37.port_b_data_in_clock = "clock1";
defparam ram_block3a37.port_b_data_out_clear = "none";
defparam ram_block3a37.port_b_data_out_clock = "none";
defparam ram_block3a37.port_b_data_width = 1;
defparam ram_block3a37.port_b_first_address = 0;
defparam ram_block3a37.port_b_first_bit_number = 5;
defparam ram_block3a37.port_b_last_address = 8191;
defparam ram_block3a37.port_b_logical_ram_depth = 16384;
defparam ram_block3a37.port_b_logical_ram_width = 32;
defparam ram_block3a37.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_read_enable_clock = "clock1";
defparam ram_block3a37.port_b_write_enable_clock = "clock1";
defparam ram_block3a37.ram_block_type = "M9K";
defparam ram_block3a37.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y33_N0
cycloneive_ram_block ram_block3a5(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a5_PORTADATAOUT_bus),
	.portbdataout(ram_block3a5_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a5.clk0_core_clock_enable = "ena0";
defparam ram_block3a5.clk1_core_clock_enable = "ena1";
defparam ram_block3a5.data_interleave_offset_in_bits = 1;
defparam ram_block3a5.data_interleave_width_in_bits = 1;
defparam ram_block3a5.init_file = "meminit.hex";
defparam ram_block3a5.init_file_layout = "port_a";
defparam ram_block3a5.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a5.operation_mode = "bidir_dual_port";
defparam ram_block3a5.port_a_address_clear = "none";
defparam ram_block3a5.port_a_address_width = 13;
defparam ram_block3a5.port_a_byte_enable_clock = "none";
defparam ram_block3a5.port_a_data_out_clear = "none";
defparam ram_block3a5.port_a_data_out_clock = "none";
defparam ram_block3a5.port_a_data_width = 1;
defparam ram_block3a5.port_a_first_address = 0;
defparam ram_block3a5.port_a_first_bit_number = 5;
defparam ram_block3a5.port_a_last_address = 8191;
defparam ram_block3a5.port_a_logical_ram_depth = 16384;
defparam ram_block3a5.port_a_logical_ram_width = 32;
defparam ram_block3a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_address_clear = "none";
defparam ram_block3a5.port_b_address_clock = "clock1";
defparam ram_block3a5.port_b_address_width = 13;
defparam ram_block3a5.port_b_data_in_clock = "clock1";
defparam ram_block3a5.port_b_data_out_clear = "none";
defparam ram_block3a5.port_b_data_out_clock = "none";
defparam ram_block3a5.port_b_data_width = 1;
defparam ram_block3a5.port_b_first_address = 0;
defparam ram_block3a5.port_b_first_bit_number = 5;
defparam ram_block3a5.port_b_last_address = 8191;
defparam ram_block3a5.port_b_logical_ram_depth = 16384;
defparam ram_block3a5.port_b_logical_ram_width = 32;
defparam ram_block3a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_read_enable_clock = "clock1";
defparam ram_block3a5.port_b_write_enable_clock = "clock1";
defparam ram_block3a5.ram_block_type = "M9K";
defparam ram_block3a5.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001C010EBB;
// synopsys translate_on

// Location: M9K_X51_Y45_N0
cycloneive_ram_block ram_block3a38(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a38_PORTADATAOUT_bus),
	.portbdataout(ram_block3a38_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a38.clk0_core_clock_enable = "ena0";
defparam ram_block3a38.clk1_core_clock_enable = "ena1";
defparam ram_block3a38.data_interleave_offset_in_bits = 1;
defparam ram_block3a38.data_interleave_width_in_bits = 1;
defparam ram_block3a38.init_file = "meminit.hex";
defparam ram_block3a38.init_file_layout = "port_a";
defparam ram_block3a38.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a38.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a38.operation_mode = "bidir_dual_port";
defparam ram_block3a38.port_a_address_clear = "none";
defparam ram_block3a38.port_a_address_width = 13;
defparam ram_block3a38.port_a_byte_enable_clock = "none";
defparam ram_block3a38.port_a_data_out_clear = "none";
defparam ram_block3a38.port_a_data_out_clock = "none";
defparam ram_block3a38.port_a_data_width = 1;
defparam ram_block3a38.port_a_first_address = 0;
defparam ram_block3a38.port_a_first_bit_number = 6;
defparam ram_block3a38.port_a_last_address = 8191;
defparam ram_block3a38.port_a_logical_ram_depth = 16384;
defparam ram_block3a38.port_a_logical_ram_width = 32;
defparam ram_block3a38.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_address_clear = "none";
defparam ram_block3a38.port_b_address_clock = "clock1";
defparam ram_block3a38.port_b_address_width = 13;
defparam ram_block3a38.port_b_data_in_clock = "clock1";
defparam ram_block3a38.port_b_data_out_clear = "none";
defparam ram_block3a38.port_b_data_out_clock = "none";
defparam ram_block3a38.port_b_data_width = 1;
defparam ram_block3a38.port_b_first_address = 0;
defparam ram_block3a38.port_b_first_bit_number = 6;
defparam ram_block3a38.port_b_last_address = 8191;
defparam ram_block3a38.port_b_logical_ram_depth = 16384;
defparam ram_block3a38.port_b_logical_ram_width = 32;
defparam ram_block3a38.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_read_enable_clock = "clock1";
defparam ram_block3a38.port_b_write_enable_clock = "clock1";
defparam ram_block3a38.ram_block_type = "M9K";
defparam ram_block3a38.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y38_N0
cycloneive_ram_block ram_block3a6(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a6_PORTADATAOUT_bus),
	.portbdataout(ram_block3a6_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a6.clk0_core_clock_enable = "ena0";
defparam ram_block3a6.clk1_core_clock_enable = "ena1";
defparam ram_block3a6.data_interleave_offset_in_bits = 1;
defparam ram_block3a6.data_interleave_width_in_bits = 1;
defparam ram_block3a6.init_file = "meminit.hex";
defparam ram_block3a6.init_file_layout = "port_a";
defparam ram_block3a6.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a6.operation_mode = "bidir_dual_port";
defparam ram_block3a6.port_a_address_clear = "none";
defparam ram_block3a6.port_a_address_width = 13;
defparam ram_block3a6.port_a_byte_enable_clock = "none";
defparam ram_block3a6.port_a_data_out_clear = "none";
defparam ram_block3a6.port_a_data_out_clock = "none";
defparam ram_block3a6.port_a_data_width = 1;
defparam ram_block3a6.port_a_first_address = 0;
defparam ram_block3a6.port_a_first_bit_number = 6;
defparam ram_block3a6.port_a_last_address = 8191;
defparam ram_block3a6.port_a_logical_ram_depth = 16384;
defparam ram_block3a6.port_a_logical_ram_width = 32;
defparam ram_block3a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_address_clear = "none";
defparam ram_block3a6.port_b_address_clock = "clock1";
defparam ram_block3a6.port_b_address_width = 13;
defparam ram_block3a6.port_b_data_in_clock = "clock1";
defparam ram_block3a6.port_b_data_out_clear = "none";
defparam ram_block3a6.port_b_data_out_clock = "none";
defparam ram_block3a6.port_b_data_width = 1;
defparam ram_block3a6.port_b_first_address = 0;
defparam ram_block3a6.port_b_first_bit_number = 6;
defparam ram_block3a6.port_b_last_address = 8191;
defparam ram_block3a6.port_b_logical_ram_depth = 16384;
defparam ram_block3a6.port_b_logical_ram_width = 32;
defparam ram_block3a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_read_enable_clock = "clock1";
defparam ram_block3a6.port_b_write_enable_clock = "clock1";
defparam ram_block3a6.ram_block_type = "M9K";
defparam ram_block3a6.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010B;
// synopsys translate_on

// Location: M9K_X51_Y43_N0
cycloneive_ram_block ram_block3a39(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a39_PORTADATAOUT_bus),
	.portbdataout(ram_block3a39_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a39.clk0_core_clock_enable = "ena0";
defparam ram_block3a39.clk1_core_clock_enable = "ena1";
defparam ram_block3a39.data_interleave_offset_in_bits = 1;
defparam ram_block3a39.data_interleave_width_in_bits = 1;
defparam ram_block3a39.init_file = "meminit.hex";
defparam ram_block3a39.init_file_layout = "port_a";
defparam ram_block3a39.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a39.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a39.operation_mode = "bidir_dual_port";
defparam ram_block3a39.port_a_address_clear = "none";
defparam ram_block3a39.port_a_address_width = 13;
defparam ram_block3a39.port_a_byte_enable_clock = "none";
defparam ram_block3a39.port_a_data_out_clear = "none";
defparam ram_block3a39.port_a_data_out_clock = "none";
defparam ram_block3a39.port_a_data_width = 1;
defparam ram_block3a39.port_a_first_address = 0;
defparam ram_block3a39.port_a_first_bit_number = 7;
defparam ram_block3a39.port_a_last_address = 8191;
defparam ram_block3a39.port_a_logical_ram_depth = 16384;
defparam ram_block3a39.port_a_logical_ram_width = 32;
defparam ram_block3a39.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_address_clear = "none";
defparam ram_block3a39.port_b_address_clock = "clock1";
defparam ram_block3a39.port_b_address_width = 13;
defparam ram_block3a39.port_b_data_in_clock = "clock1";
defparam ram_block3a39.port_b_data_out_clear = "none";
defparam ram_block3a39.port_b_data_out_clock = "none";
defparam ram_block3a39.port_b_data_width = 1;
defparam ram_block3a39.port_b_first_address = 0;
defparam ram_block3a39.port_b_first_bit_number = 7;
defparam ram_block3a39.port_b_last_address = 8191;
defparam ram_block3a39.port_b_logical_ram_depth = 16384;
defparam ram_block3a39.port_b_logical_ram_width = 32;
defparam ram_block3a39.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_read_enable_clock = "clock1";
defparam ram_block3a39.port_b_write_enable_clock = "clock1";
defparam ram_block3a39.ram_block_type = "M9K";
defparam ram_block3a39.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y44_N0
cycloneive_ram_block ram_block3a7(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a7_PORTADATAOUT_bus),
	.portbdataout(ram_block3a7_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a7.clk0_core_clock_enable = "ena0";
defparam ram_block3a7.clk1_core_clock_enable = "ena1";
defparam ram_block3a7.data_interleave_offset_in_bits = 1;
defparam ram_block3a7.data_interleave_width_in_bits = 1;
defparam ram_block3a7.init_file = "meminit.hex";
defparam ram_block3a7.init_file_layout = "port_a";
defparam ram_block3a7.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a7.operation_mode = "bidir_dual_port";
defparam ram_block3a7.port_a_address_clear = "none";
defparam ram_block3a7.port_a_address_width = 13;
defparam ram_block3a7.port_a_byte_enable_clock = "none";
defparam ram_block3a7.port_a_data_out_clear = "none";
defparam ram_block3a7.port_a_data_out_clock = "none";
defparam ram_block3a7.port_a_data_width = 1;
defparam ram_block3a7.port_a_first_address = 0;
defparam ram_block3a7.port_a_first_bit_number = 7;
defparam ram_block3a7.port_a_last_address = 8191;
defparam ram_block3a7.port_a_logical_ram_depth = 16384;
defparam ram_block3a7.port_a_logical_ram_width = 32;
defparam ram_block3a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_address_clear = "none";
defparam ram_block3a7.port_b_address_clock = "clock1";
defparam ram_block3a7.port_b_address_width = 13;
defparam ram_block3a7.port_b_data_in_clock = "clock1";
defparam ram_block3a7.port_b_data_out_clear = "none";
defparam ram_block3a7.port_b_data_out_clock = "none";
defparam ram_block3a7.port_b_data_width = 1;
defparam ram_block3a7.port_b_first_address = 0;
defparam ram_block3a7.port_b_first_bit_number = 7;
defparam ram_block3a7.port_b_last_address = 8191;
defparam ram_block3a7.port_b_logical_ram_depth = 16384;
defparam ram_block3a7.port_b_logical_ram_width = 32;
defparam ram_block3a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_read_enable_clock = "clock1";
defparam ram_block3a7.port_b_write_enable_clock = "clock1";
defparam ram_block3a7.ram_block_type = "M9K";
defparam ram_block3a7.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000E;
// synopsys translate_on

// Location: M9K_X51_Y47_N0
cycloneive_ram_block ram_block3a40(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a40_PORTADATAOUT_bus),
	.portbdataout(ram_block3a40_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a40.clk0_core_clock_enable = "ena0";
defparam ram_block3a40.clk1_core_clock_enable = "ena1";
defparam ram_block3a40.data_interleave_offset_in_bits = 1;
defparam ram_block3a40.data_interleave_width_in_bits = 1;
defparam ram_block3a40.init_file = "meminit.hex";
defparam ram_block3a40.init_file_layout = "port_a";
defparam ram_block3a40.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a40.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a40.operation_mode = "bidir_dual_port";
defparam ram_block3a40.port_a_address_clear = "none";
defparam ram_block3a40.port_a_address_width = 13;
defparam ram_block3a40.port_a_byte_enable_clock = "none";
defparam ram_block3a40.port_a_data_out_clear = "none";
defparam ram_block3a40.port_a_data_out_clock = "none";
defparam ram_block3a40.port_a_data_width = 1;
defparam ram_block3a40.port_a_first_address = 0;
defparam ram_block3a40.port_a_first_bit_number = 8;
defparam ram_block3a40.port_a_last_address = 8191;
defparam ram_block3a40.port_a_logical_ram_depth = 16384;
defparam ram_block3a40.port_a_logical_ram_width = 32;
defparam ram_block3a40.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_address_clear = "none";
defparam ram_block3a40.port_b_address_clock = "clock1";
defparam ram_block3a40.port_b_address_width = 13;
defparam ram_block3a40.port_b_data_in_clock = "clock1";
defparam ram_block3a40.port_b_data_out_clear = "none";
defparam ram_block3a40.port_b_data_out_clock = "none";
defparam ram_block3a40.port_b_data_width = 1;
defparam ram_block3a40.port_b_first_address = 0;
defparam ram_block3a40.port_b_first_bit_number = 8;
defparam ram_block3a40.port_b_last_address = 8191;
defparam ram_block3a40.port_b_logical_ram_depth = 16384;
defparam ram_block3a40.port_b_logical_ram_width = 32;
defparam ram_block3a40.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_read_enable_clock = "clock1";
defparam ram_block3a40.port_b_write_enable_clock = "clock1";
defparam ram_block3a40.ram_block_type = "M9K";
defparam ram_block3a40.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y36_N0
cycloneive_ram_block ram_block3a8(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a8_PORTADATAOUT_bus),
	.portbdataout(ram_block3a8_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a8.clk0_core_clock_enable = "ena0";
defparam ram_block3a8.clk1_core_clock_enable = "ena1";
defparam ram_block3a8.data_interleave_offset_in_bits = 1;
defparam ram_block3a8.data_interleave_width_in_bits = 1;
defparam ram_block3a8.init_file = "meminit.hex";
defparam ram_block3a8.init_file_layout = "port_a";
defparam ram_block3a8.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a8.operation_mode = "bidir_dual_port";
defparam ram_block3a8.port_a_address_clear = "none";
defparam ram_block3a8.port_a_address_width = 13;
defparam ram_block3a8.port_a_byte_enable_clock = "none";
defparam ram_block3a8.port_a_data_out_clear = "none";
defparam ram_block3a8.port_a_data_out_clock = "none";
defparam ram_block3a8.port_a_data_width = 1;
defparam ram_block3a8.port_a_first_address = 0;
defparam ram_block3a8.port_a_first_bit_number = 8;
defparam ram_block3a8.port_a_last_address = 8191;
defparam ram_block3a8.port_a_logical_ram_depth = 16384;
defparam ram_block3a8.port_a_logical_ram_width = 32;
defparam ram_block3a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_address_clear = "none";
defparam ram_block3a8.port_b_address_clock = "clock1";
defparam ram_block3a8.port_b_address_width = 13;
defparam ram_block3a8.port_b_data_in_clock = "clock1";
defparam ram_block3a8.port_b_data_out_clear = "none";
defparam ram_block3a8.port_b_data_out_clock = "none";
defparam ram_block3a8.port_b_data_width = 1;
defparam ram_block3a8.port_b_first_address = 0;
defparam ram_block3a8.port_b_first_bit_number = 8;
defparam ram_block3a8.port_b_last_address = 8191;
defparam ram_block3a8.port_b_logical_ram_depth = 16384;
defparam ram_block3a8.port_b_logical_ram_width = 32;
defparam ram_block3a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_read_enable_clock = "clock1";
defparam ram_block3a8.port_b_write_enable_clock = "clock1";
defparam ram_block3a8.ram_block_type = "M9K";
defparam ram_block3a8.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000902;
// synopsys translate_on

// Location: M9K_X51_Y39_N0
cycloneive_ram_block ram_block3a41(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a41_PORTADATAOUT_bus),
	.portbdataout(ram_block3a41_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a41.clk0_core_clock_enable = "ena0";
defparam ram_block3a41.clk1_core_clock_enable = "ena1";
defparam ram_block3a41.data_interleave_offset_in_bits = 1;
defparam ram_block3a41.data_interleave_width_in_bits = 1;
defparam ram_block3a41.init_file = "meminit.hex";
defparam ram_block3a41.init_file_layout = "port_a";
defparam ram_block3a41.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a41.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a41.operation_mode = "bidir_dual_port";
defparam ram_block3a41.port_a_address_clear = "none";
defparam ram_block3a41.port_a_address_width = 13;
defparam ram_block3a41.port_a_byte_enable_clock = "none";
defparam ram_block3a41.port_a_data_out_clear = "none";
defparam ram_block3a41.port_a_data_out_clock = "none";
defparam ram_block3a41.port_a_data_width = 1;
defparam ram_block3a41.port_a_first_address = 0;
defparam ram_block3a41.port_a_first_bit_number = 9;
defparam ram_block3a41.port_a_last_address = 8191;
defparam ram_block3a41.port_a_logical_ram_depth = 16384;
defparam ram_block3a41.port_a_logical_ram_width = 32;
defparam ram_block3a41.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_address_clear = "none";
defparam ram_block3a41.port_b_address_clock = "clock1";
defparam ram_block3a41.port_b_address_width = 13;
defparam ram_block3a41.port_b_data_in_clock = "clock1";
defparam ram_block3a41.port_b_data_out_clear = "none";
defparam ram_block3a41.port_b_data_out_clock = "none";
defparam ram_block3a41.port_b_data_width = 1;
defparam ram_block3a41.port_b_first_address = 0;
defparam ram_block3a41.port_b_first_bit_number = 9;
defparam ram_block3a41.port_b_last_address = 8191;
defparam ram_block3a41.port_b_logical_ram_depth = 16384;
defparam ram_block3a41.port_b_logical_ram_width = 32;
defparam ram_block3a41.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_read_enable_clock = "clock1";
defparam ram_block3a41.port_b_write_enable_clock = "clock1";
defparam ram_block3a41.ram_block_type = "M9K";
defparam ram_block3a41.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y33_N0
cycloneive_ram_block ram_block3a9(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a9_PORTADATAOUT_bus),
	.portbdataout(ram_block3a9_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a9.clk0_core_clock_enable = "ena0";
defparam ram_block3a9.clk1_core_clock_enable = "ena1";
defparam ram_block3a9.data_interleave_offset_in_bits = 1;
defparam ram_block3a9.data_interleave_width_in_bits = 1;
defparam ram_block3a9.init_file = "meminit.hex";
defparam ram_block3a9.init_file_layout = "port_a";
defparam ram_block3a9.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a9.operation_mode = "bidir_dual_port";
defparam ram_block3a9.port_a_address_clear = "none";
defparam ram_block3a9.port_a_address_width = 13;
defparam ram_block3a9.port_a_byte_enable_clock = "none";
defparam ram_block3a9.port_a_data_out_clear = "none";
defparam ram_block3a9.port_a_data_out_clock = "none";
defparam ram_block3a9.port_a_data_width = 1;
defparam ram_block3a9.port_a_first_address = 0;
defparam ram_block3a9.port_a_first_bit_number = 9;
defparam ram_block3a9.port_a_last_address = 8191;
defparam ram_block3a9.port_a_logical_ram_depth = 16384;
defparam ram_block3a9.port_a_logical_ram_width = 32;
defparam ram_block3a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_address_clear = "none";
defparam ram_block3a9.port_b_address_clock = "clock1";
defparam ram_block3a9.port_b_address_width = 13;
defparam ram_block3a9.port_b_data_in_clock = "clock1";
defparam ram_block3a9.port_b_data_out_clear = "none";
defparam ram_block3a9.port_b_data_out_clock = "none";
defparam ram_block3a9.port_b_data_width = 1;
defparam ram_block3a9.port_b_first_address = 0;
defparam ram_block3a9.port_b_first_bit_number = 9;
defparam ram_block3a9.port_b_last_address = 8191;
defparam ram_block3a9.port_b_logical_ram_depth = 16384;
defparam ram_block3a9.port_b_logical_ram_width = 32;
defparam ram_block3a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_read_enable_clock = "clock1";
defparam ram_block3a9.port_b_write_enable_clock = "clock1";
defparam ram_block3a9.ram_block_type = "M9K";
defparam ram_block3a9.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000903;
// synopsys translate_on

// Location: M9K_X37_Y37_N0
cycloneive_ram_block ram_block3a42(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a42_PORTADATAOUT_bus),
	.portbdataout(ram_block3a42_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a42.clk0_core_clock_enable = "ena0";
defparam ram_block3a42.clk1_core_clock_enable = "ena1";
defparam ram_block3a42.data_interleave_offset_in_bits = 1;
defparam ram_block3a42.data_interleave_width_in_bits = 1;
defparam ram_block3a42.init_file = "meminit.hex";
defparam ram_block3a42.init_file_layout = "port_a";
defparam ram_block3a42.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a42.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a42.operation_mode = "bidir_dual_port";
defparam ram_block3a42.port_a_address_clear = "none";
defparam ram_block3a42.port_a_address_width = 13;
defparam ram_block3a42.port_a_byte_enable_clock = "none";
defparam ram_block3a42.port_a_data_out_clear = "none";
defparam ram_block3a42.port_a_data_out_clock = "none";
defparam ram_block3a42.port_a_data_width = 1;
defparam ram_block3a42.port_a_first_address = 0;
defparam ram_block3a42.port_a_first_bit_number = 10;
defparam ram_block3a42.port_a_last_address = 8191;
defparam ram_block3a42.port_a_logical_ram_depth = 16384;
defparam ram_block3a42.port_a_logical_ram_width = 32;
defparam ram_block3a42.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_address_clear = "none";
defparam ram_block3a42.port_b_address_clock = "clock1";
defparam ram_block3a42.port_b_address_width = 13;
defparam ram_block3a42.port_b_data_in_clock = "clock1";
defparam ram_block3a42.port_b_data_out_clear = "none";
defparam ram_block3a42.port_b_data_out_clock = "none";
defparam ram_block3a42.port_b_data_width = 1;
defparam ram_block3a42.port_b_first_address = 0;
defparam ram_block3a42.port_b_first_bit_number = 10;
defparam ram_block3a42.port_b_last_address = 8191;
defparam ram_block3a42.port_b_logical_ram_depth = 16384;
defparam ram_block3a42.port_b_logical_ram_width = 32;
defparam ram_block3a42.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_read_enable_clock = "clock1";
defparam ram_block3a42.port_b_write_enable_clock = "clock1";
defparam ram_block3a42.ram_block_type = "M9K";
defparam ram_block3a42.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y41_N0
cycloneive_ram_block ram_block3a10(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a10_PORTADATAOUT_bus),
	.portbdataout(ram_block3a10_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a10.clk0_core_clock_enable = "ena0";
defparam ram_block3a10.clk1_core_clock_enable = "ena1";
defparam ram_block3a10.data_interleave_offset_in_bits = 1;
defparam ram_block3a10.data_interleave_width_in_bits = 1;
defparam ram_block3a10.init_file = "meminit.hex";
defparam ram_block3a10.init_file_layout = "port_a";
defparam ram_block3a10.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a10.operation_mode = "bidir_dual_port";
defparam ram_block3a10.port_a_address_clear = "none";
defparam ram_block3a10.port_a_address_width = 13;
defparam ram_block3a10.port_a_byte_enable_clock = "none";
defparam ram_block3a10.port_a_data_out_clear = "none";
defparam ram_block3a10.port_a_data_out_clock = "none";
defparam ram_block3a10.port_a_data_width = 1;
defparam ram_block3a10.port_a_first_address = 0;
defparam ram_block3a10.port_a_first_bit_number = 10;
defparam ram_block3a10.port_a_last_address = 8191;
defparam ram_block3a10.port_a_logical_ram_depth = 16384;
defparam ram_block3a10.port_a_logical_ram_width = 32;
defparam ram_block3a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_address_clear = "none";
defparam ram_block3a10.port_b_address_clock = "clock1";
defparam ram_block3a10.port_b_address_width = 13;
defparam ram_block3a10.port_b_data_in_clock = "clock1";
defparam ram_block3a10.port_b_data_out_clear = "none";
defparam ram_block3a10.port_b_data_out_clock = "none";
defparam ram_block3a10.port_b_data_width = 1;
defparam ram_block3a10.port_b_first_address = 0;
defparam ram_block3a10.port_b_first_bit_number = 10;
defparam ram_block3a10.port_b_last_address = 8191;
defparam ram_block3a10.port_b_logical_ram_depth = 16384;
defparam ram_block3a10.port_b_logical_ram_width = 32;
defparam ram_block3a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_read_enable_clock = "clock1";
defparam ram_block3a10.port_b_write_enable_clock = "clock1";
defparam ram_block3a10.ram_block_type = "M9K";
defparam ram_block3a10.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000102;
// synopsys translate_on

// Location: M9K_X51_Y49_N0
cycloneive_ram_block ram_block3a43(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a43_PORTADATAOUT_bus),
	.portbdataout(ram_block3a43_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a43.clk0_core_clock_enable = "ena0";
defparam ram_block3a43.clk1_core_clock_enable = "ena1";
defparam ram_block3a43.data_interleave_offset_in_bits = 1;
defparam ram_block3a43.data_interleave_width_in_bits = 1;
defparam ram_block3a43.init_file = "meminit.hex";
defparam ram_block3a43.init_file_layout = "port_a";
defparam ram_block3a43.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a43.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a43.operation_mode = "bidir_dual_port";
defparam ram_block3a43.port_a_address_clear = "none";
defparam ram_block3a43.port_a_address_width = 13;
defparam ram_block3a43.port_a_byte_enable_clock = "none";
defparam ram_block3a43.port_a_data_out_clear = "none";
defparam ram_block3a43.port_a_data_out_clock = "none";
defparam ram_block3a43.port_a_data_width = 1;
defparam ram_block3a43.port_a_first_address = 0;
defparam ram_block3a43.port_a_first_bit_number = 11;
defparam ram_block3a43.port_a_last_address = 8191;
defparam ram_block3a43.port_a_logical_ram_depth = 16384;
defparam ram_block3a43.port_a_logical_ram_width = 32;
defparam ram_block3a43.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_address_clear = "none";
defparam ram_block3a43.port_b_address_clock = "clock1";
defparam ram_block3a43.port_b_address_width = 13;
defparam ram_block3a43.port_b_data_in_clock = "clock1";
defparam ram_block3a43.port_b_data_out_clear = "none";
defparam ram_block3a43.port_b_data_out_clock = "none";
defparam ram_block3a43.port_b_data_width = 1;
defparam ram_block3a43.port_b_first_address = 0;
defparam ram_block3a43.port_b_first_bit_number = 11;
defparam ram_block3a43.port_b_last_address = 8191;
defparam ram_block3a43.port_b_logical_ram_depth = 16384;
defparam ram_block3a43.port_b_logical_ram_width = 32;
defparam ram_block3a43.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_read_enable_clock = "clock1";
defparam ram_block3a43.port_b_write_enable_clock = "clock1";
defparam ram_block3a43.ram_block_type = "M9K";
defparam ram_block3a43.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y48_N0
cycloneive_ram_block ram_block3a11(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a11_PORTADATAOUT_bus),
	.portbdataout(ram_block3a11_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a11.clk0_core_clock_enable = "ena0";
defparam ram_block3a11.clk1_core_clock_enable = "ena1";
defparam ram_block3a11.data_interleave_offset_in_bits = 1;
defparam ram_block3a11.data_interleave_width_in_bits = 1;
defparam ram_block3a11.init_file = "meminit.hex";
defparam ram_block3a11.init_file_layout = "port_a";
defparam ram_block3a11.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a11.operation_mode = "bidir_dual_port";
defparam ram_block3a11.port_a_address_clear = "none";
defparam ram_block3a11.port_a_address_width = 13;
defparam ram_block3a11.port_a_byte_enable_clock = "none";
defparam ram_block3a11.port_a_data_out_clear = "none";
defparam ram_block3a11.port_a_data_out_clock = "none";
defparam ram_block3a11.port_a_data_width = 1;
defparam ram_block3a11.port_a_first_address = 0;
defparam ram_block3a11.port_a_first_bit_number = 11;
defparam ram_block3a11.port_a_last_address = 8191;
defparam ram_block3a11.port_a_logical_ram_depth = 16384;
defparam ram_block3a11.port_a_logical_ram_width = 32;
defparam ram_block3a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_address_clear = "none";
defparam ram_block3a11.port_b_address_clock = "clock1";
defparam ram_block3a11.port_b_address_width = 13;
defparam ram_block3a11.port_b_data_in_clock = "clock1";
defparam ram_block3a11.port_b_data_out_clear = "none";
defparam ram_block3a11.port_b_data_out_clock = "none";
defparam ram_block3a11.port_b_data_width = 1;
defparam ram_block3a11.port_b_first_address = 0;
defparam ram_block3a11.port_b_first_bit_number = 11;
defparam ram_block3a11.port_b_last_address = 8191;
defparam ram_block3a11.port_b_logical_ram_depth = 16384;
defparam ram_block3a11.port_b_logical_ram_width = 32;
defparam ram_block3a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_read_enable_clock = "clock1";
defparam ram_block3a11.port_b_write_enable_clock = "clock1";
defparam ram_block3a11.ram_block_type = "M9K";
defparam ram_block3a11.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010012410;
// synopsys translate_on

// Location: M9K_X64_Y41_N0
cycloneive_ram_block ram_block3a44(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a44_PORTADATAOUT_bus),
	.portbdataout(ram_block3a44_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a44.clk0_core_clock_enable = "ena0";
defparam ram_block3a44.clk1_core_clock_enable = "ena1";
defparam ram_block3a44.data_interleave_offset_in_bits = 1;
defparam ram_block3a44.data_interleave_width_in_bits = 1;
defparam ram_block3a44.init_file = "meminit.hex";
defparam ram_block3a44.init_file_layout = "port_a";
defparam ram_block3a44.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a44.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a44.operation_mode = "bidir_dual_port";
defparam ram_block3a44.port_a_address_clear = "none";
defparam ram_block3a44.port_a_address_width = 13;
defparam ram_block3a44.port_a_byte_enable_clock = "none";
defparam ram_block3a44.port_a_data_out_clear = "none";
defparam ram_block3a44.port_a_data_out_clock = "none";
defparam ram_block3a44.port_a_data_width = 1;
defparam ram_block3a44.port_a_first_address = 0;
defparam ram_block3a44.port_a_first_bit_number = 12;
defparam ram_block3a44.port_a_last_address = 8191;
defparam ram_block3a44.port_a_logical_ram_depth = 16384;
defparam ram_block3a44.port_a_logical_ram_width = 32;
defparam ram_block3a44.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_address_clear = "none";
defparam ram_block3a44.port_b_address_clock = "clock1";
defparam ram_block3a44.port_b_address_width = 13;
defparam ram_block3a44.port_b_data_in_clock = "clock1";
defparam ram_block3a44.port_b_data_out_clear = "none";
defparam ram_block3a44.port_b_data_out_clock = "none";
defparam ram_block3a44.port_b_data_width = 1;
defparam ram_block3a44.port_b_first_address = 0;
defparam ram_block3a44.port_b_first_bit_number = 12;
defparam ram_block3a44.port_b_last_address = 8191;
defparam ram_block3a44.port_b_logical_ram_depth = 16384;
defparam ram_block3a44.port_b_logical_ram_width = 32;
defparam ram_block3a44.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_read_enable_clock = "clock1";
defparam ram_block3a44.port_b_write_enable_clock = "clock1";
defparam ram_block3a44.ram_block_type = "M9K";
defparam ram_block3a44.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y39_N0
cycloneive_ram_block ram_block3a12(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a12_PORTADATAOUT_bus),
	.portbdataout(ram_block3a12_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a12.clk0_core_clock_enable = "ena0";
defparam ram_block3a12.clk1_core_clock_enable = "ena1";
defparam ram_block3a12.data_interleave_offset_in_bits = 1;
defparam ram_block3a12.data_interleave_width_in_bits = 1;
defparam ram_block3a12.init_file = "meminit.hex";
defparam ram_block3a12.init_file_layout = "port_a";
defparam ram_block3a12.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a12.operation_mode = "bidir_dual_port";
defparam ram_block3a12.port_a_address_clear = "none";
defparam ram_block3a12.port_a_address_width = 13;
defparam ram_block3a12.port_a_byte_enable_clock = "none";
defparam ram_block3a12.port_a_data_out_clear = "none";
defparam ram_block3a12.port_a_data_out_clock = "none";
defparam ram_block3a12.port_a_data_width = 1;
defparam ram_block3a12.port_a_first_address = 0;
defparam ram_block3a12.port_a_first_bit_number = 12;
defparam ram_block3a12.port_a_last_address = 8191;
defparam ram_block3a12.port_a_logical_ram_depth = 16384;
defparam ram_block3a12.port_a_logical_ram_width = 32;
defparam ram_block3a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_address_clear = "none";
defparam ram_block3a12.port_b_address_clock = "clock1";
defparam ram_block3a12.port_b_address_width = 13;
defparam ram_block3a12.port_b_data_in_clock = "clock1";
defparam ram_block3a12.port_b_data_out_clear = "none";
defparam ram_block3a12.port_b_data_out_clock = "none";
defparam ram_block3a12.port_b_data_width = 1;
defparam ram_block3a12.port_b_first_address = 0;
defparam ram_block3a12.port_b_first_bit_number = 12;
defparam ram_block3a12.port_b_last_address = 8191;
defparam ram_block3a12.port_b_logical_ram_depth = 16384;
defparam ram_block3a12.port_b_logical_ram_width = 32;
defparam ram_block3a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_read_enable_clock = "clock1";
defparam ram_block3a12.port_b_write_enable_clock = "clock1";
defparam ram_block3a12.ram_block_type = "M9K";
defparam ram_block3a12.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010002893;
// synopsys translate_on

// Location: M9K_X64_Y35_N0
cycloneive_ram_block ram_block3a45(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a45_PORTADATAOUT_bus),
	.portbdataout(ram_block3a45_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a45.clk0_core_clock_enable = "ena0";
defparam ram_block3a45.clk1_core_clock_enable = "ena1";
defparam ram_block3a45.data_interleave_offset_in_bits = 1;
defparam ram_block3a45.data_interleave_width_in_bits = 1;
defparam ram_block3a45.init_file = "meminit.hex";
defparam ram_block3a45.init_file_layout = "port_a";
defparam ram_block3a45.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a45.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a45.operation_mode = "bidir_dual_port";
defparam ram_block3a45.port_a_address_clear = "none";
defparam ram_block3a45.port_a_address_width = 13;
defparam ram_block3a45.port_a_byte_enable_clock = "none";
defparam ram_block3a45.port_a_data_out_clear = "none";
defparam ram_block3a45.port_a_data_out_clock = "none";
defparam ram_block3a45.port_a_data_width = 1;
defparam ram_block3a45.port_a_first_address = 0;
defparam ram_block3a45.port_a_first_bit_number = 13;
defparam ram_block3a45.port_a_last_address = 8191;
defparam ram_block3a45.port_a_logical_ram_depth = 16384;
defparam ram_block3a45.port_a_logical_ram_width = 32;
defparam ram_block3a45.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_address_clear = "none";
defparam ram_block3a45.port_b_address_clock = "clock1";
defparam ram_block3a45.port_b_address_width = 13;
defparam ram_block3a45.port_b_data_in_clock = "clock1";
defparam ram_block3a45.port_b_data_out_clear = "none";
defparam ram_block3a45.port_b_data_out_clock = "none";
defparam ram_block3a45.port_b_data_width = 1;
defparam ram_block3a45.port_b_first_address = 0;
defparam ram_block3a45.port_b_first_bit_number = 13;
defparam ram_block3a45.port_b_last_address = 8191;
defparam ram_block3a45.port_b_logical_ram_depth = 16384;
defparam ram_block3a45.port_b_logical_ram_width = 32;
defparam ram_block3a45.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_read_enable_clock = "clock1";
defparam ram_block3a45.port_b_write_enable_clock = "clock1";
defparam ram_block3a45.ram_block_type = "M9K";
defparam ram_block3a45.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y45_N0
cycloneive_ram_block ram_block3a13(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a13_PORTADATAOUT_bus),
	.portbdataout(ram_block3a13_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a13.clk0_core_clock_enable = "ena0";
defparam ram_block3a13.clk1_core_clock_enable = "ena1";
defparam ram_block3a13.data_interleave_offset_in_bits = 1;
defparam ram_block3a13.data_interleave_width_in_bits = 1;
defparam ram_block3a13.init_file = "meminit.hex";
defparam ram_block3a13.init_file_layout = "port_a";
defparam ram_block3a13.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a13.operation_mode = "bidir_dual_port";
defparam ram_block3a13.port_a_address_clear = "none";
defparam ram_block3a13.port_a_address_width = 13;
defparam ram_block3a13.port_a_byte_enable_clock = "none";
defparam ram_block3a13.port_a_data_out_clear = "none";
defparam ram_block3a13.port_a_data_out_clock = "none";
defparam ram_block3a13.port_a_data_width = 1;
defparam ram_block3a13.port_a_first_address = 0;
defparam ram_block3a13.port_a_first_bit_number = 13;
defparam ram_block3a13.port_a_last_address = 8191;
defparam ram_block3a13.port_a_logical_ram_depth = 16384;
defparam ram_block3a13.port_a_logical_ram_width = 32;
defparam ram_block3a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_address_clear = "none";
defparam ram_block3a13.port_b_address_clock = "clock1";
defparam ram_block3a13.port_b_address_width = 13;
defparam ram_block3a13.port_b_data_in_clock = "clock1";
defparam ram_block3a13.port_b_data_out_clear = "none";
defparam ram_block3a13.port_b_data_out_clock = "none";
defparam ram_block3a13.port_b_data_width = 1;
defparam ram_block3a13.port_b_first_address = 0;
defparam ram_block3a13.port_b_first_bit_number = 13;
defparam ram_block3a13.port_b_last_address = 8191;
defparam ram_block3a13.port_b_logical_ram_depth = 16384;
defparam ram_block3a13.port_b_logical_ram_width = 32;
defparam ram_block3a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_read_enable_clock = "clock1";
defparam ram_block3a13.port_b_write_enable_clock = "clock1";
defparam ram_block3a13.ram_block_type = "M9K";
defparam ram_block3a13.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100188A2;
// synopsys translate_on

// Location: M9K_X51_Y27_N0
cycloneive_ram_block ram_block3a46(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a46_PORTADATAOUT_bus),
	.portbdataout(ram_block3a46_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a46.clk0_core_clock_enable = "ena0";
defparam ram_block3a46.clk1_core_clock_enable = "ena1";
defparam ram_block3a46.data_interleave_offset_in_bits = 1;
defparam ram_block3a46.data_interleave_width_in_bits = 1;
defparam ram_block3a46.init_file = "meminit.hex";
defparam ram_block3a46.init_file_layout = "port_a";
defparam ram_block3a46.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a46.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a46.operation_mode = "bidir_dual_port";
defparam ram_block3a46.port_a_address_clear = "none";
defparam ram_block3a46.port_a_address_width = 13;
defparam ram_block3a46.port_a_byte_enable_clock = "none";
defparam ram_block3a46.port_a_data_out_clear = "none";
defparam ram_block3a46.port_a_data_out_clock = "none";
defparam ram_block3a46.port_a_data_width = 1;
defparam ram_block3a46.port_a_first_address = 0;
defparam ram_block3a46.port_a_first_bit_number = 14;
defparam ram_block3a46.port_a_last_address = 8191;
defparam ram_block3a46.port_a_logical_ram_depth = 16384;
defparam ram_block3a46.port_a_logical_ram_width = 32;
defparam ram_block3a46.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_address_clear = "none";
defparam ram_block3a46.port_b_address_clock = "clock1";
defparam ram_block3a46.port_b_address_width = 13;
defparam ram_block3a46.port_b_data_in_clock = "clock1";
defparam ram_block3a46.port_b_data_out_clear = "none";
defparam ram_block3a46.port_b_data_out_clock = "none";
defparam ram_block3a46.port_b_data_width = 1;
defparam ram_block3a46.port_b_first_address = 0;
defparam ram_block3a46.port_b_first_bit_number = 14;
defparam ram_block3a46.port_b_last_address = 8191;
defparam ram_block3a46.port_b_logical_ram_depth = 16384;
defparam ram_block3a46.port_b_logical_ram_width = 32;
defparam ram_block3a46.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_read_enable_clock = "clock1";
defparam ram_block3a46.port_b_write_enable_clock = "clock1";
defparam ram_block3a46.ram_block_type = "M9K";
defparam ram_block3a46.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y28_N0
cycloneive_ram_block ram_block3a14(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a14_PORTADATAOUT_bus),
	.portbdataout(ram_block3a14_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a14.clk0_core_clock_enable = "ena0";
defparam ram_block3a14.clk1_core_clock_enable = "ena1";
defparam ram_block3a14.data_interleave_offset_in_bits = 1;
defparam ram_block3a14.data_interleave_width_in_bits = 1;
defparam ram_block3a14.init_file = "meminit.hex";
defparam ram_block3a14.init_file_layout = "port_a";
defparam ram_block3a14.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a14.operation_mode = "bidir_dual_port";
defparam ram_block3a14.port_a_address_clear = "none";
defparam ram_block3a14.port_a_address_width = 13;
defparam ram_block3a14.port_a_byte_enable_clock = "none";
defparam ram_block3a14.port_a_data_out_clear = "none";
defparam ram_block3a14.port_a_data_out_clock = "none";
defparam ram_block3a14.port_a_data_width = 1;
defparam ram_block3a14.port_a_first_address = 0;
defparam ram_block3a14.port_a_first_bit_number = 14;
defparam ram_block3a14.port_a_last_address = 8191;
defparam ram_block3a14.port_a_logical_ram_depth = 16384;
defparam ram_block3a14.port_a_logical_ram_width = 32;
defparam ram_block3a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_address_clear = "none";
defparam ram_block3a14.port_b_address_clock = "clock1";
defparam ram_block3a14.port_b_address_width = 13;
defparam ram_block3a14.port_b_data_in_clock = "clock1";
defparam ram_block3a14.port_b_data_out_clear = "none";
defparam ram_block3a14.port_b_data_out_clock = "none";
defparam ram_block3a14.port_b_data_width = 1;
defparam ram_block3a14.port_b_first_address = 0;
defparam ram_block3a14.port_b_first_bit_number = 14;
defparam ram_block3a14.port_b_last_address = 8191;
defparam ram_block3a14.port_b_logical_ram_depth = 16384;
defparam ram_block3a14.port_b_logical_ram_width = 32;
defparam ram_block3a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_read_enable_clock = "clock1";
defparam ram_block3a14.port_b_write_enable_clock = "clock1";
defparam ram_block3a14.ram_block_type = "M9K";
defparam ram_block3a14.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001AE01;
// synopsys translate_on

// Location: M9K_X78_Y30_N0
cycloneive_ram_block ram_block3a47(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a47_PORTADATAOUT_bus),
	.portbdataout(ram_block3a47_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a47.clk0_core_clock_enable = "ena0";
defparam ram_block3a47.clk1_core_clock_enable = "ena1";
defparam ram_block3a47.data_interleave_offset_in_bits = 1;
defparam ram_block3a47.data_interleave_width_in_bits = 1;
defparam ram_block3a47.init_file = "meminit.hex";
defparam ram_block3a47.init_file_layout = "port_a";
defparam ram_block3a47.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a47.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a47.operation_mode = "bidir_dual_port";
defparam ram_block3a47.port_a_address_clear = "none";
defparam ram_block3a47.port_a_address_width = 13;
defparam ram_block3a47.port_a_byte_enable_clock = "none";
defparam ram_block3a47.port_a_data_out_clear = "none";
defparam ram_block3a47.port_a_data_out_clock = "none";
defparam ram_block3a47.port_a_data_width = 1;
defparam ram_block3a47.port_a_first_address = 0;
defparam ram_block3a47.port_a_first_bit_number = 15;
defparam ram_block3a47.port_a_last_address = 8191;
defparam ram_block3a47.port_a_logical_ram_depth = 16384;
defparam ram_block3a47.port_a_logical_ram_width = 32;
defparam ram_block3a47.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_address_clear = "none";
defparam ram_block3a47.port_b_address_clock = "clock1";
defparam ram_block3a47.port_b_address_width = 13;
defparam ram_block3a47.port_b_data_in_clock = "clock1";
defparam ram_block3a47.port_b_data_out_clear = "none";
defparam ram_block3a47.port_b_data_out_clock = "none";
defparam ram_block3a47.port_b_data_width = 1;
defparam ram_block3a47.port_b_first_address = 0;
defparam ram_block3a47.port_b_first_bit_number = 15;
defparam ram_block3a47.port_b_last_address = 8191;
defparam ram_block3a47.port_b_logical_ram_depth = 16384;
defparam ram_block3a47.port_b_logical_ram_width = 32;
defparam ram_block3a47.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_read_enable_clock = "clock1";
defparam ram_block3a47.port_b_write_enable_clock = "clock1";
defparam ram_block3a47.ram_block_type = "M9K";
defparam ram_block3a47.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y28_N0
cycloneive_ram_block ram_block3a15(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a15_PORTADATAOUT_bus),
	.portbdataout(ram_block3a15_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a15.clk0_core_clock_enable = "ena0";
defparam ram_block3a15.clk1_core_clock_enable = "ena1";
defparam ram_block3a15.data_interleave_offset_in_bits = 1;
defparam ram_block3a15.data_interleave_width_in_bits = 1;
defparam ram_block3a15.init_file = "meminit.hex";
defparam ram_block3a15.init_file_layout = "port_a";
defparam ram_block3a15.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a15.operation_mode = "bidir_dual_port";
defparam ram_block3a15.port_a_address_clear = "none";
defparam ram_block3a15.port_a_address_width = 13;
defparam ram_block3a15.port_a_byte_enable_clock = "none";
defparam ram_block3a15.port_a_data_out_clear = "none";
defparam ram_block3a15.port_a_data_out_clock = "none";
defparam ram_block3a15.port_a_data_width = 1;
defparam ram_block3a15.port_a_first_address = 0;
defparam ram_block3a15.port_a_first_bit_number = 15;
defparam ram_block3a15.port_a_last_address = 8191;
defparam ram_block3a15.port_a_logical_ram_depth = 16384;
defparam ram_block3a15.port_a_logical_ram_width = 32;
defparam ram_block3a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_address_clear = "none";
defparam ram_block3a15.port_b_address_clock = "clock1";
defparam ram_block3a15.port_b_address_width = 13;
defparam ram_block3a15.port_b_data_in_clock = "clock1";
defparam ram_block3a15.port_b_data_out_clear = "none";
defparam ram_block3a15.port_b_data_out_clock = "none";
defparam ram_block3a15.port_b_data_width = 1;
defparam ram_block3a15.port_b_first_address = 0;
defparam ram_block3a15.port_b_first_bit_number = 15;
defparam ram_block3a15.port_b_last_address = 8191;
defparam ram_block3a15.port_b_logical_ram_depth = 16384;
defparam ram_block3a15.port_b_logical_ram_width = 32;
defparam ram_block3a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_read_enable_clock = "clock1";
defparam ram_block3a15.port_b_write_enable_clock = "clock1";
defparam ram_block3a15.ram_block_type = "M9K";
defparam ram_block3a15.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000901;
// synopsys translate_on

// Location: M9K_X51_Y32_N0
cycloneive_ram_block ram_block3a48(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a48_PORTADATAOUT_bus),
	.portbdataout(ram_block3a48_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a48.clk0_core_clock_enable = "ena0";
defparam ram_block3a48.clk1_core_clock_enable = "ena1";
defparam ram_block3a48.data_interleave_offset_in_bits = 1;
defparam ram_block3a48.data_interleave_width_in_bits = 1;
defparam ram_block3a48.init_file = "meminit.hex";
defparam ram_block3a48.init_file_layout = "port_a";
defparam ram_block3a48.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a48.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a48.operation_mode = "bidir_dual_port";
defparam ram_block3a48.port_a_address_clear = "none";
defparam ram_block3a48.port_a_address_width = 13;
defparam ram_block3a48.port_a_byte_enable_clock = "none";
defparam ram_block3a48.port_a_data_out_clear = "none";
defparam ram_block3a48.port_a_data_out_clock = "none";
defparam ram_block3a48.port_a_data_width = 1;
defparam ram_block3a48.port_a_first_address = 0;
defparam ram_block3a48.port_a_first_bit_number = 16;
defparam ram_block3a48.port_a_last_address = 8191;
defparam ram_block3a48.port_a_logical_ram_depth = 16384;
defparam ram_block3a48.port_a_logical_ram_width = 32;
defparam ram_block3a48.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_address_clear = "none";
defparam ram_block3a48.port_b_address_clock = "clock1";
defparam ram_block3a48.port_b_address_width = 13;
defparam ram_block3a48.port_b_data_in_clock = "clock1";
defparam ram_block3a48.port_b_data_out_clear = "none";
defparam ram_block3a48.port_b_data_out_clock = "none";
defparam ram_block3a48.port_b_data_width = 1;
defparam ram_block3a48.port_b_first_address = 0;
defparam ram_block3a48.port_b_first_bit_number = 16;
defparam ram_block3a48.port_b_last_address = 8191;
defparam ram_block3a48.port_b_logical_ram_depth = 16384;
defparam ram_block3a48.port_b_logical_ram_width = 32;
defparam ram_block3a48.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_read_enable_clock = "clock1";
defparam ram_block3a48.port_b_write_enable_clock = "clock1";
defparam ram_block3a48.ram_block_type = "M9K";
defparam ram_block3a48.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y30_N0
cycloneive_ram_block ram_block3a16(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a16_PORTADATAOUT_bus),
	.portbdataout(ram_block3a16_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a16.clk0_core_clock_enable = "ena0";
defparam ram_block3a16.clk1_core_clock_enable = "ena1";
defparam ram_block3a16.data_interleave_offset_in_bits = 1;
defparam ram_block3a16.data_interleave_width_in_bits = 1;
defparam ram_block3a16.init_file = "meminit.hex";
defparam ram_block3a16.init_file_layout = "port_a";
defparam ram_block3a16.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a16.operation_mode = "bidir_dual_port";
defparam ram_block3a16.port_a_address_clear = "none";
defparam ram_block3a16.port_a_address_width = 13;
defparam ram_block3a16.port_a_byte_enable_clock = "none";
defparam ram_block3a16.port_a_data_out_clear = "none";
defparam ram_block3a16.port_a_data_out_clock = "none";
defparam ram_block3a16.port_a_data_width = 1;
defparam ram_block3a16.port_a_first_address = 0;
defparam ram_block3a16.port_a_first_bit_number = 16;
defparam ram_block3a16.port_a_last_address = 8191;
defparam ram_block3a16.port_a_logical_ram_depth = 16384;
defparam ram_block3a16.port_a_logical_ram_width = 32;
defparam ram_block3a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_address_clear = "none";
defparam ram_block3a16.port_b_address_clock = "clock1";
defparam ram_block3a16.port_b_address_width = 13;
defparam ram_block3a16.port_b_data_in_clock = "clock1";
defparam ram_block3a16.port_b_data_out_clear = "none";
defparam ram_block3a16.port_b_data_out_clock = "none";
defparam ram_block3a16.port_b_data_width = 1;
defparam ram_block3a16.port_b_first_address = 0;
defparam ram_block3a16.port_b_first_bit_number = 16;
defparam ram_block3a16.port_b_last_address = 8191;
defparam ram_block3a16.port_b_logical_ram_depth = 16384;
defparam ram_block3a16.port_b_logical_ram_width = 32;
defparam ram_block3a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_read_enable_clock = "clock1";
defparam ram_block3a16.port_b_write_enable_clock = "clock1";
defparam ram_block3a16.ram_block_type = "M9K";
defparam ram_block3a16.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001556A145;
// synopsys translate_on

// Location: M9K_X64_Y31_N0
cycloneive_ram_block ram_block3a49(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a49_PORTADATAOUT_bus),
	.portbdataout(ram_block3a49_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a49.clk0_core_clock_enable = "ena0";
defparam ram_block3a49.clk1_core_clock_enable = "ena1";
defparam ram_block3a49.data_interleave_offset_in_bits = 1;
defparam ram_block3a49.data_interleave_width_in_bits = 1;
defparam ram_block3a49.init_file = "meminit.hex";
defparam ram_block3a49.init_file_layout = "port_a";
defparam ram_block3a49.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a49.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a49.operation_mode = "bidir_dual_port";
defparam ram_block3a49.port_a_address_clear = "none";
defparam ram_block3a49.port_a_address_width = 13;
defparam ram_block3a49.port_a_byte_enable_clock = "none";
defparam ram_block3a49.port_a_data_out_clear = "none";
defparam ram_block3a49.port_a_data_out_clock = "none";
defparam ram_block3a49.port_a_data_width = 1;
defparam ram_block3a49.port_a_first_address = 0;
defparam ram_block3a49.port_a_first_bit_number = 17;
defparam ram_block3a49.port_a_last_address = 8191;
defparam ram_block3a49.port_a_logical_ram_depth = 16384;
defparam ram_block3a49.port_a_logical_ram_width = 32;
defparam ram_block3a49.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_address_clear = "none";
defparam ram_block3a49.port_b_address_clock = "clock1";
defparam ram_block3a49.port_b_address_width = 13;
defparam ram_block3a49.port_b_data_in_clock = "clock1";
defparam ram_block3a49.port_b_data_out_clear = "none";
defparam ram_block3a49.port_b_data_out_clock = "none";
defparam ram_block3a49.port_b_data_width = 1;
defparam ram_block3a49.port_b_first_address = 0;
defparam ram_block3a49.port_b_first_bit_number = 17;
defparam ram_block3a49.port_b_last_address = 8191;
defparam ram_block3a49.port_b_logical_ram_depth = 16384;
defparam ram_block3a49.port_b_logical_ram_width = 32;
defparam ram_block3a49.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_read_enable_clock = "clock1";
defparam ram_block3a49.port_b_write_enable_clock = "clock1";
defparam ram_block3a49.ram_block_type = "M9K";
defparam ram_block3a49.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y34_N0
cycloneive_ram_block ram_block3a17(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a17_PORTADATAOUT_bus),
	.portbdataout(ram_block3a17_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a17.clk0_core_clock_enable = "ena0";
defparam ram_block3a17.clk1_core_clock_enable = "ena1";
defparam ram_block3a17.data_interleave_offset_in_bits = 1;
defparam ram_block3a17.data_interleave_width_in_bits = 1;
defparam ram_block3a17.init_file = "meminit.hex";
defparam ram_block3a17.init_file_layout = "port_a";
defparam ram_block3a17.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a17.operation_mode = "bidir_dual_port";
defparam ram_block3a17.port_a_address_clear = "none";
defparam ram_block3a17.port_a_address_width = 13;
defparam ram_block3a17.port_a_byte_enable_clock = "none";
defparam ram_block3a17.port_a_data_out_clear = "none";
defparam ram_block3a17.port_a_data_out_clock = "none";
defparam ram_block3a17.port_a_data_width = 1;
defparam ram_block3a17.port_a_first_address = 0;
defparam ram_block3a17.port_a_first_bit_number = 17;
defparam ram_block3a17.port_a_last_address = 8191;
defparam ram_block3a17.port_a_logical_ram_depth = 16384;
defparam ram_block3a17.port_a_logical_ram_width = 32;
defparam ram_block3a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_address_clear = "none";
defparam ram_block3a17.port_b_address_clock = "clock1";
defparam ram_block3a17.port_b_address_width = 13;
defparam ram_block3a17.port_b_data_in_clock = "clock1";
defparam ram_block3a17.port_b_data_out_clear = "none";
defparam ram_block3a17.port_b_data_out_clock = "none";
defparam ram_block3a17.port_b_data_width = 1;
defparam ram_block3a17.port_b_first_address = 0;
defparam ram_block3a17.port_b_first_bit_number = 17;
defparam ram_block3a17.port_b_last_address = 8191;
defparam ram_block3a17.port_b_logical_ram_depth = 16384;
defparam ram_block3a17.port_b_logical_ram_width = 32;
defparam ram_block3a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_read_enable_clock = "clock1";
defparam ram_block3a17.port_b_write_enable_clock = "clock1";
defparam ram_block3a17.ram_block_type = "M9K";
defparam ram_block3a17.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000016655FBA;
// synopsys translate_on

// Location: M9K_X51_Y25_N0
cycloneive_ram_block ram_block3a50(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a50_PORTADATAOUT_bus),
	.portbdataout(ram_block3a50_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a50.clk0_core_clock_enable = "ena0";
defparam ram_block3a50.clk1_core_clock_enable = "ena1";
defparam ram_block3a50.data_interleave_offset_in_bits = 1;
defparam ram_block3a50.data_interleave_width_in_bits = 1;
defparam ram_block3a50.init_file = "meminit.hex";
defparam ram_block3a50.init_file_layout = "port_a";
defparam ram_block3a50.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a50.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a50.operation_mode = "bidir_dual_port";
defparam ram_block3a50.port_a_address_clear = "none";
defparam ram_block3a50.port_a_address_width = 13;
defparam ram_block3a50.port_a_byte_enable_clock = "none";
defparam ram_block3a50.port_a_data_out_clear = "none";
defparam ram_block3a50.port_a_data_out_clock = "none";
defparam ram_block3a50.port_a_data_width = 1;
defparam ram_block3a50.port_a_first_address = 0;
defparam ram_block3a50.port_a_first_bit_number = 18;
defparam ram_block3a50.port_a_last_address = 8191;
defparam ram_block3a50.port_a_logical_ram_depth = 16384;
defparam ram_block3a50.port_a_logical_ram_width = 32;
defparam ram_block3a50.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_address_clear = "none";
defparam ram_block3a50.port_b_address_clock = "clock1";
defparam ram_block3a50.port_b_address_width = 13;
defparam ram_block3a50.port_b_data_in_clock = "clock1";
defparam ram_block3a50.port_b_data_out_clear = "none";
defparam ram_block3a50.port_b_data_out_clock = "none";
defparam ram_block3a50.port_b_data_width = 1;
defparam ram_block3a50.port_b_first_address = 0;
defparam ram_block3a50.port_b_first_bit_number = 18;
defparam ram_block3a50.port_b_last_address = 8191;
defparam ram_block3a50.port_b_logical_ram_depth = 16384;
defparam ram_block3a50.port_b_logical_ram_width = 32;
defparam ram_block3a50.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_read_enable_clock = "clock1";
defparam ram_block3a50.port_b_write_enable_clock = "clock1";
defparam ram_block3a50.ram_block_type = "M9K";
defparam ram_block3a50.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y33_N0
cycloneive_ram_block ram_block3a18(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a18_PORTADATAOUT_bus),
	.portbdataout(ram_block3a18_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a18.clk0_core_clock_enable = "ena0";
defparam ram_block3a18.clk1_core_clock_enable = "ena1";
defparam ram_block3a18.data_interleave_offset_in_bits = 1;
defparam ram_block3a18.data_interleave_width_in_bits = 1;
defparam ram_block3a18.init_file = "meminit.hex";
defparam ram_block3a18.init_file_layout = "port_a";
defparam ram_block3a18.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a18.operation_mode = "bidir_dual_port";
defparam ram_block3a18.port_a_address_clear = "none";
defparam ram_block3a18.port_a_address_width = 13;
defparam ram_block3a18.port_a_byte_enable_clock = "none";
defparam ram_block3a18.port_a_data_out_clear = "none";
defparam ram_block3a18.port_a_data_out_clock = "none";
defparam ram_block3a18.port_a_data_width = 1;
defparam ram_block3a18.port_a_first_address = 0;
defparam ram_block3a18.port_a_first_bit_number = 18;
defparam ram_block3a18.port_a_last_address = 8191;
defparam ram_block3a18.port_a_logical_ram_depth = 16384;
defparam ram_block3a18.port_a_logical_ram_width = 32;
defparam ram_block3a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_address_clear = "none";
defparam ram_block3a18.port_b_address_clock = "clock1";
defparam ram_block3a18.port_b_address_width = 13;
defparam ram_block3a18.port_b_data_in_clock = "clock1";
defparam ram_block3a18.port_b_data_out_clear = "none";
defparam ram_block3a18.port_b_data_out_clock = "none";
defparam ram_block3a18.port_b_data_width = 1;
defparam ram_block3a18.port_b_first_address = 0;
defparam ram_block3a18.port_b_first_bit_number = 18;
defparam ram_block3a18.port_b_last_address = 8191;
defparam ram_block3a18.port_b_logical_ram_depth = 16384;
defparam ram_block3a18.port_b_logical_ram_width = 32;
defparam ram_block3a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_read_enable_clock = "clock1";
defparam ram_block3a18.port_b_write_enable_clock = "clock1";
defparam ram_block3a18.ram_block_type = "M9K";
defparam ram_block3a18.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000187A514C;
// synopsys translate_on

// Location: M9K_X51_Y33_N0
cycloneive_ram_block ram_block3a51(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a51_PORTADATAOUT_bus),
	.portbdataout(ram_block3a51_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a51.clk0_core_clock_enable = "ena0";
defparam ram_block3a51.clk1_core_clock_enable = "ena1";
defparam ram_block3a51.data_interleave_offset_in_bits = 1;
defparam ram_block3a51.data_interleave_width_in_bits = 1;
defparam ram_block3a51.init_file = "meminit.hex";
defparam ram_block3a51.init_file_layout = "port_a";
defparam ram_block3a51.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a51.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a51.operation_mode = "bidir_dual_port";
defparam ram_block3a51.port_a_address_clear = "none";
defparam ram_block3a51.port_a_address_width = 13;
defparam ram_block3a51.port_a_byte_enable_clock = "none";
defparam ram_block3a51.port_a_data_out_clear = "none";
defparam ram_block3a51.port_a_data_out_clock = "none";
defparam ram_block3a51.port_a_data_width = 1;
defparam ram_block3a51.port_a_first_address = 0;
defparam ram_block3a51.port_a_first_bit_number = 19;
defparam ram_block3a51.port_a_last_address = 8191;
defparam ram_block3a51.port_a_logical_ram_depth = 16384;
defparam ram_block3a51.port_a_logical_ram_width = 32;
defparam ram_block3a51.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_address_clear = "none";
defparam ram_block3a51.port_b_address_clock = "clock1";
defparam ram_block3a51.port_b_address_width = 13;
defparam ram_block3a51.port_b_data_in_clock = "clock1";
defparam ram_block3a51.port_b_data_out_clear = "none";
defparam ram_block3a51.port_b_data_out_clock = "none";
defparam ram_block3a51.port_b_data_width = 1;
defparam ram_block3a51.port_b_first_address = 0;
defparam ram_block3a51.port_b_first_bit_number = 19;
defparam ram_block3a51.port_b_last_address = 8191;
defparam ram_block3a51.port_b_logical_ram_depth = 16384;
defparam ram_block3a51.port_b_logical_ram_width = 32;
defparam ram_block3a51.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_read_enable_clock = "clock1";
defparam ram_block3a51.port_b_write_enable_clock = "clock1";
defparam ram_block3a51.ram_block_type = "M9K";
defparam ram_block3a51.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y35_N0
cycloneive_ram_block ram_block3a19(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a19_PORTADATAOUT_bus),
	.portbdataout(ram_block3a19_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a19.clk0_core_clock_enable = "ena0";
defparam ram_block3a19.clk1_core_clock_enable = "ena1";
defparam ram_block3a19.data_interleave_offset_in_bits = 1;
defparam ram_block3a19.data_interleave_width_in_bits = 1;
defparam ram_block3a19.init_file = "meminit.hex";
defparam ram_block3a19.init_file_layout = "port_a";
defparam ram_block3a19.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a19.operation_mode = "bidir_dual_port";
defparam ram_block3a19.port_a_address_clear = "none";
defparam ram_block3a19.port_a_address_width = 13;
defparam ram_block3a19.port_a_byte_enable_clock = "none";
defparam ram_block3a19.port_a_data_out_clear = "none";
defparam ram_block3a19.port_a_data_out_clock = "none";
defparam ram_block3a19.port_a_data_width = 1;
defparam ram_block3a19.port_a_first_address = 0;
defparam ram_block3a19.port_a_first_bit_number = 19;
defparam ram_block3a19.port_a_last_address = 8191;
defparam ram_block3a19.port_a_logical_ram_depth = 16384;
defparam ram_block3a19.port_a_logical_ram_width = 32;
defparam ram_block3a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_address_clear = "none";
defparam ram_block3a19.port_b_address_clock = "clock1";
defparam ram_block3a19.port_b_address_width = 13;
defparam ram_block3a19.port_b_data_in_clock = "clock1";
defparam ram_block3a19.port_b_data_out_clear = "none";
defparam ram_block3a19.port_b_data_out_clock = "none";
defparam ram_block3a19.port_b_data_width = 1;
defparam ram_block3a19.port_b_first_address = 0;
defparam ram_block3a19.port_b_first_bit_number = 19;
defparam ram_block3a19.port_b_last_address = 8191;
defparam ram_block3a19.port_b_logical_ram_depth = 16384;
defparam ram_block3a19.port_b_logical_ram_width = 32;
defparam ram_block3a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_read_enable_clock = "clock1";
defparam ram_block3a19.port_b_write_enable_clock = "clock1";
defparam ram_block3a19.ram_block_type = "M9K";
defparam ram_block3a19.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001F825800;
// synopsys translate_on

// Location: M9K_X37_Y31_N0
cycloneive_ram_block ram_block3a52(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a52_PORTADATAOUT_bus),
	.portbdataout(ram_block3a52_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a52.clk0_core_clock_enable = "ena0";
defparam ram_block3a52.clk1_core_clock_enable = "ena1";
defparam ram_block3a52.data_interleave_offset_in_bits = 1;
defparam ram_block3a52.data_interleave_width_in_bits = 1;
defparam ram_block3a52.init_file = "meminit.hex";
defparam ram_block3a52.init_file_layout = "port_a";
defparam ram_block3a52.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a52.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a52.operation_mode = "bidir_dual_port";
defparam ram_block3a52.port_a_address_clear = "none";
defparam ram_block3a52.port_a_address_width = 13;
defparam ram_block3a52.port_a_byte_enable_clock = "none";
defparam ram_block3a52.port_a_data_out_clear = "none";
defparam ram_block3a52.port_a_data_out_clock = "none";
defparam ram_block3a52.port_a_data_width = 1;
defparam ram_block3a52.port_a_first_address = 0;
defparam ram_block3a52.port_a_first_bit_number = 20;
defparam ram_block3a52.port_a_last_address = 8191;
defparam ram_block3a52.port_a_logical_ram_depth = 16384;
defparam ram_block3a52.port_a_logical_ram_width = 32;
defparam ram_block3a52.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_address_clear = "none";
defparam ram_block3a52.port_b_address_clock = "clock1";
defparam ram_block3a52.port_b_address_width = 13;
defparam ram_block3a52.port_b_data_in_clock = "clock1";
defparam ram_block3a52.port_b_data_out_clear = "none";
defparam ram_block3a52.port_b_data_out_clock = "none";
defparam ram_block3a52.port_b_data_width = 1;
defparam ram_block3a52.port_b_first_address = 0;
defparam ram_block3a52.port_b_first_bit_number = 20;
defparam ram_block3a52.port_b_last_address = 8191;
defparam ram_block3a52.port_b_logical_ram_depth = 16384;
defparam ram_block3a52.port_b_logical_ram_width = 32;
defparam ram_block3a52.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_read_enable_clock = "clock1";
defparam ram_block3a52.port_b_write_enable_clock = "clock1";
defparam ram_block3a52.ram_block_type = "M9K";
defparam ram_block3a52.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y31_N0
cycloneive_ram_block ram_block3a20(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a20_PORTADATAOUT_bus),
	.portbdataout(ram_block3a20_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a20.clk0_core_clock_enable = "ena0";
defparam ram_block3a20.clk1_core_clock_enable = "ena1";
defparam ram_block3a20.data_interleave_offset_in_bits = 1;
defparam ram_block3a20.data_interleave_width_in_bits = 1;
defparam ram_block3a20.init_file = "meminit.hex";
defparam ram_block3a20.init_file_layout = "port_a";
defparam ram_block3a20.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a20.operation_mode = "bidir_dual_port";
defparam ram_block3a20.port_a_address_clear = "none";
defparam ram_block3a20.port_a_address_width = 13;
defparam ram_block3a20.port_a_byte_enable_clock = "none";
defparam ram_block3a20.port_a_data_out_clear = "none";
defparam ram_block3a20.port_a_data_out_clock = "none";
defparam ram_block3a20.port_a_data_width = 1;
defparam ram_block3a20.port_a_first_address = 0;
defparam ram_block3a20.port_a_first_bit_number = 20;
defparam ram_block3a20.port_a_last_address = 8191;
defparam ram_block3a20.port_a_logical_ram_depth = 16384;
defparam ram_block3a20.port_a_logical_ram_width = 32;
defparam ram_block3a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_address_clear = "none";
defparam ram_block3a20.port_b_address_clock = "clock1";
defparam ram_block3a20.port_b_address_width = 13;
defparam ram_block3a20.port_b_data_in_clock = "clock1";
defparam ram_block3a20.port_b_data_out_clear = "none";
defparam ram_block3a20.port_b_data_out_clock = "none";
defparam ram_block3a20.port_b_data_width = 1;
defparam ram_block3a20.port_b_first_address = 0;
defparam ram_block3a20.port_b_first_bit_number = 20;
defparam ram_block3a20.port_b_last_address = 8191;
defparam ram_block3a20.port_b_logical_ram_depth = 16384;
defparam ram_block3a20.port_b_logical_ram_width = 32;
defparam ram_block3a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_read_enable_clock = "clock1";
defparam ram_block3a20.port_b_write_enable_clock = "clock1";
defparam ram_block3a20.ram_block_type = "M9K";
defparam ram_block3a20.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000C;
// synopsys translate_on

// Location: M9K_X51_Y37_N0
cycloneive_ram_block ram_block3a53(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a53_PORTADATAOUT_bus),
	.portbdataout(ram_block3a53_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a53.clk0_core_clock_enable = "ena0";
defparam ram_block3a53.clk1_core_clock_enable = "ena1";
defparam ram_block3a53.data_interleave_offset_in_bits = 1;
defparam ram_block3a53.data_interleave_width_in_bits = 1;
defparam ram_block3a53.init_file = "meminit.hex";
defparam ram_block3a53.init_file_layout = "port_a";
defparam ram_block3a53.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a53.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a53.operation_mode = "bidir_dual_port";
defparam ram_block3a53.port_a_address_clear = "none";
defparam ram_block3a53.port_a_address_width = 13;
defparam ram_block3a53.port_a_byte_enable_clock = "none";
defparam ram_block3a53.port_a_data_out_clear = "none";
defparam ram_block3a53.port_a_data_out_clock = "none";
defparam ram_block3a53.port_a_data_width = 1;
defparam ram_block3a53.port_a_first_address = 0;
defparam ram_block3a53.port_a_first_bit_number = 21;
defparam ram_block3a53.port_a_last_address = 8191;
defparam ram_block3a53.port_a_logical_ram_depth = 16384;
defparam ram_block3a53.port_a_logical_ram_width = 32;
defparam ram_block3a53.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_address_clear = "none";
defparam ram_block3a53.port_b_address_clock = "clock1";
defparam ram_block3a53.port_b_address_width = 13;
defparam ram_block3a53.port_b_data_in_clock = "clock1";
defparam ram_block3a53.port_b_data_out_clear = "none";
defparam ram_block3a53.port_b_data_out_clock = "none";
defparam ram_block3a53.port_b_data_width = 1;
defparam ram_block3a53.port_b_first_address = 0;
defparam ram_block3a53.port_b_first_bit_number = 21;
defparam ram_block3a53.port_b_last_address = 8191;
defparam ram_block3a53.port_b_logical_ram_depth = 16384;
defparam ram_block3a53.port_b_logical_ram_width = 32;
defparam ram_block3a53.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_read_enable_clock = "clock1";
defparam ram_block3a53.port_b_write_enable_clock = "clock1";
defparam ram_block3a53.ram_block_type = "M9K";
defparam ram_block3a53.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y37_N0
cycloneive_ram_block ram_block3a21(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a21_PORTADATAOUT_bus),
	.portbdataout(ram_block3a21_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a21.clk0_core_clock_enable = "ena0";
defparam ram_block3a21.clk1_core_clock_enable = "ena1";
defparam ram_block3a21.data_interleave_offset_in_bits = 1;
defparam ram_block3a21.data_interleave_width_in_bits = 1;
defparam ram_block3a21.init_file = "meminit.hex";
defparam ram_block3a21.init_file_layout = "port_a";
defparam ram_block3a21.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a21.operation_mode = "bidir_dual_port";
defparam ram_block3a21.port_a_address_clear = "none";
defparam ram_block3a21.port_a_address_width = 13;
defparam ram_block3a21.port_a_byte_enable_clock = "none";
defparam ram_block3a21.port_a_data_out_clear = "none";
defparam ram_block3a21.port_a_data_out_clock = "none";
defparam ram_block3a21.port_a_data_width = 1;
defparam ram_block3a21.port_a_first_address = 0;
defparam ram_block3a21.port_a_first_bit_number = 21;
defparam ram_block3a21.port_a_last_address = 8191;
defparam ram_block3a21.port_a_logical_ram_depth = 16384;
defparam ram_block3a21.port_a_logical_ram_width = 32;
defparam ram_block3a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_address_clear = "none";
defparam ram_block3a21.port_b_address_clock = "clock1";
defparam ram_block3a21.port_b_address_width = 13;
defparam ram_block3a21.port_b_data_in_clock = "clock1";
defparam ram_block3a21.port_b_data_out_clear = "none";
defparam ram_block3a21.port_b_data_out_clock = "none";
defparam ram_block3a21.port_b_data_width = 1;
defparam ram_block3a21.port_b_first_address = 0;
defparam ram_block3a21.port_b_first_bit_number = 21;
defparam ram_block3a21.port_b_last_address = 8191;
defparam ram_block3a21.port_b_logical_ram_depth = 16384;
defparam ram_block3a21.port_b_logical_ram_width = 32;
defparam ram_block3a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_read_enable_clock = "clock1";
defparam ram_block3a21.port_b_write_enable_clock = "clock1";
defparam ram_block3a21.ram_block_type = "M9K";
defparam ram_block3a21.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFD0DF0;
// synopsys translate_on

// Location: M9K_X51_Y36_N0
cycloneive_ram_block ram_block3a54(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a54_PORTADATAOUT_bus),
	.portbdataout(ram_block3a54_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a54.clk0_core_clock_enable = "ena0";
defparam ram_block3a54.clk1_core_clock_enable = "ena1";
defparam ram_block3a54.data_interleave_offset_in_bits = 1;
defparam ram_block3a54.data_interleave_width_in_bits = 1;
defparam ram_block3a54.init_file = "meminit.hex";
defparam ram_block3a54.init_file_layout = "port_a";
defparam ram_block3a54.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a54.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a54.operation_mode = "bidir_dual_port";
defparam ram_block3a54.port_a_address_clear = "none";
defparam ram_block3a54.port_a_address_width = 13;
defparam ram_block3a54.port_a_byte_enable_clock = "none";
defparam ram_block3a54.port_a_data_out_clear = "none";
defparam ram_block3a54.port_a_data_out_clock = "none";
defparam ram_block3a54.port_a_data_width = 1;
defparam ram_block3a54.port_a_first_address = 0;
defparam ram_block3a54.port_a_first_bit_number = 22;
defparam ram_block3a54.port_a_last_address = 8191;
defparam ram_block3a54.port_a_logical_ram_depth = 16384;
defparam ram_block3a54.port_a_logical_ram_width = 32;
defparam ram_block3a54.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_address_clear = "none";
defparam ram_block3a54.port_b_address_clock = "clock1";
defparam ram_block3a54.port_b_address_width = 13;
defparam ram_block3a54.port_b_data_in_clock = "clock1";
defparam ram_block3a54.port_b_data_out_clear = "none";
defparam ram_block3a54.port_b_data_out_clock = "none";
defparam ram_block3a54.port_b_data_width = 1;
defparam ram_block3a54.port_b_first_address = 0;
defparam ram_block3a54.port_b_first_bit_number = 22;
defparam ram_block3a54.port_b_last_address = 8191;
defparam ram_block3a54.port_b_logical_ram_depth = 16384;
defparam ram_block3a54.port_b_logical_ram_width = 32;
defparam ram_block3a54.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_read_enable_clock = "clock1";
defparam ram_block3a54.port_b_write_enable_clock = "clock1";
defparam ram_block3a54.ram_block_type = "M9K";
defparam ram_block3a54.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y36_N0
cycloneive_ram_block ram_block3a22(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a22_PORTADATAOUT_bus),
	.portbdataout(ram_block3a22_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a22.clk0_core_clock_enable = "ena0";
defparam ram_block3a22.clk1_core_clock_enable = "ena1";
defparam ram_block3a22.data_interleave_offset_in_bits = 1;
defparam ram_block3a22.data_interleave_width_in_bits = 1;
defparam ram_block3a22.init_file = "meminit.hex";
defparam ram_block3a22.init_file_layout = "port_a";
defparam ram_block3a22.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a22.operation_mode = "bidir_dual_port";
defparam ram_block3a22.port_a_address_clear = "none";
defparam ram_block3a22.port_a_address_width = 13;
defparam ram_block3a22.port_a_byte_enable_clock = "none";
defparam ram_block3a22.port_a_data_out_clear = "none";
defparam ram_block3a22.port_a_data_out_clock = "none";
defparam ram_block3a22.port_a_data_width = 1;
defparam ram_block3a22.port_a_first_address = 0;
defparam ram_block3a22.port_a_first_bit_number = 22;
defparam ram_block3a22.port_a_last_address = 8191;
defparam ram_block3a22.port_a_logical_ram_depth = 16384;
defparam ram_block3a22.port_a_logical_ram_width = 32;
defparam ram_block3a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_address_clear = "none";
defparam ram_block3a22.port_b_address_clock = "clock1";
defparam ram_block3a22.port_b_address_width = 13;
defparam ram_block3a22.port_b_data_in_clock = "clock1";
defparam ram_block3a22.port_b_data_out_clear = "none";
defparam ram_block3a22.port_b_data_out_clock = "none";
defparam ram_block3a22.port_b_data_width = 1;
defparam ram_block3a22.port_b_first_address = 0;
defparam ram_block3a22.port_b_first_bit_number = 22;
defparam ram_block3a22.port_b_last_address = 8191;
defparam ram_block3a22.port_b_logical_ram_depth = 16384;
defparam ram_block3a22.port_b_logical_ram_width = 32;
defparam ram_block3a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_read_enable_clock = "clock1";
defparam ram_block3a22.port_b_write_enable_clock = "clock1";
defparam ram_block3a22.ram_block_type = "M9K";
defparam ram_block3a22.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001002A100;
// synopsys translate_on

// Location: M9K_X78_Y37_N0
cycloneive_ram_block ram_block3a55(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a55_PORTADATAOUT_bus),
	.portbdataout(ram_block3a55_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a55.clk0_core_clock_enable = "ena0";
defparam ram_block3a55.clk1_core_clock_enable = "ena1";
defparam ram_block3a55.data_interleave_offset_in_bits = 1;
defparam ram_block3a55.data_interleave_width_in_bits = 1;
defparam ram_block3a55.init_file = "meminit.hex";
defparam ram_block3a55.init_file_layout = "port_a";
defparam ram_block3a55.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a55.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a55.operation_mode = "bidir_dual_port";
defparam ram_block3a55.port_a_address_clear = "none";
defparam ram_block3a55.port_a_address_width = 13;
defparam ram_block3a55.port_a_byte_enable_clock = "none";
defparam ram_block3a55.port_a_data_out_clear = "none";
defparam ram_block3a55.port_a_data_out_clock = "none";
defparam ram_block3a55.port_a_data_width = 1;
defparam ram_block3a55.port_a_first_address = 0;
defparam ram_block3a55.port_a_first_bit_number = 23;
defparam ram_block3a55.port_a_last_address = 8191;
defparam ram_block3a55.port_a_logical_ram_depth = 16384;
defparam ram_block3a55.port_a_logical_ram_width = 32;
defparam ram_block3a55.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_address_clear = "none";
defparam ram_block3a55.port_b_address_clock = "clock1";
defparam ram_block3a55.port_b_address_width = 13;
defparam ram_block3a55.port_b_data_in_clock = "clock1";
defparam ram_block3a55.port_b_data_out_clear = "none";
defparam ram_block3a55.port_b_data_out_clock = "none";
defparam ram_block3a55.port_b_data_width = 1;
defparam ram_block3a55.port_b_first_address = 0;
defparam ram_block3a55.port_b_first_bit_number = 23;
defparam ram_block3a55.port_b_last_address = 8191;
defparam ram_block3a55.port_b_logical_ram_depth = 16384;
defparam ram_block3a55.port_b_logical_ram_width = 32;
defparam ram_block3a55.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_read_enable_clock = "clock1";
defparam ram_block3a55.port_b_write_enable_clock = "clock1";
defparam ram_block3a55.ram_block_type = "M9K";
defparam ram_block3a55.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y38_N0
cycloneive_ram_block ram_block3a23(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a23_PORTADATAOUT_bus),
	.portbdataout(ram_block3a23_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a23.clk0_core_clock_enable = "ena0";
defparam ram_block3a23.clk1_core_clock_enable = "ena1";
defparam ram_block3a23.data_interleave_offset_in_bits = 1;
defparam ram_block3a23.data_interleave_width_in_bits = 1;
defparam ram_block3a23.init_file = "meminit.hex";
defparam ram_block3a23.init_file_layout = "port_a";
defparam ram_block3a23.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a23.operation_mode = "bidir_dual_port";
defparam ram_block3a23.port_a_address_clear = "none";
defparam ram_block3a23.port_a_address_width = 13;
defparam ram_block3a23.port_a_byte_enable_clock = "none";
defparam ram_block3a23.port_a_data_out_clear = "none";
defparam ram_block3a23.port_a_data_out_clock = "none";
defparam ram_block3a23.port_a_data_width = 1;
defparam ram_block3a23.port_a_first_address = 0;
defparam ram_block3a23.port_a_first_bit_number = 23;
defparam ram_block3a23.port_a_last_address = 8191;
defparam ram_block3a23.port_a_logical_ram_depth = 16384;
defparam ram_block3a23.port_a_logical_ram_width = 32;
defparam ram_block3a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_address_clear = "none";
defparam ram_block3a23.port_b_address_clock = "clock1";
defparam ram_block3a23.port_b_address_width = 13;
defparam ram_block3a23.port_b_data_in_clock = "clock1";
defparam ram_block3a23.port_b_data_out_clear = "none";
defparam ram_block3a23.port_b_data_out_clock = "none";
defparam ram_block3a23.port_b_data_width = 1;
defparam ram_block3a23.port_b_first_address = 0;
defparam ram_block3a23.port_b_first_bit_number = 23;
defparam ram_block3a23.port_b_last_address = 8191;
defparam ram_block3a23.port_b_logical_ram_depth = 16384;
defparam ram_block3a23.port_b_logical_ram_width = 32;
defparam ram_block3a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_read_enable_clock = "clock1";
defparam ram_block3a23.port_b_write_enable_clock = "clock1";
defparam ram_block3a23.ram_block_type = "M9K";
defparam ram_block3a23.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFEA600;
// synopsys translate_on

// Location: M9K_X51_Y42_N0
cycloneive_ram_block ram_block3a56(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a56_PORTADATAOUT_bus),
	.portbdataout(ram_block3a56_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a56.clk0_core_clock_enable = "ena0";
defparam ram_block3a56.clk1_core_clock_enable = "ena1";
defparam ram_block3a56.data_interleave_offset_in_bits = 1;
defparam ram_block3a56.data_interleave_width_in_bits = 1;
defparam ram_block3a56.init_file = "meminit.hex";
defparam ram_block3a56.init_file_layout = "port_a";
defparam ram_block3a56.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a56.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a56.operation_mode = "bidir_dual_port";
defparam ram_block3a56.port_a_address_clear = "none";
defparam ram_block3a56.port_a_address_width = 13;
defparam ram_block3a56.port_a_byte_enable_clock = "none";
defparam ram_block3a56.port_a_data_out_clear = "none";
defparam ram_block3a56.port_a_data_out_clock = "none";
defparam ram_block3a56.port_a_data_width = 1;
defparam ram_block3a56.port_a_first_address = 0;
defparam ram_block3a56.port_a_first_bit_number = 24;
defparam ram_block3a56.port_a_last_address = 8191;
defparam ram_block3a56.port_a_logical_ram_depth = 16384;
defparam ram_block3a56.port_a_logical_ram_width = 32;
defparam ram_block3a56.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_address_clear = "none";
defparam ram_block3a56.port_b_address_clock = "clock1";
defparam ram_block3a56.port_b_address_width = 13;
defparam ram_block3a56.port_b_data_in_clock = "clock1";
defparam ram_block3a56.port_b_data_out_clear = "none";
defparam ram_block3a56.port_b_data_out_clock = "none";
defparam ram_block3a56.port_b_data_width = 1;
defparam ram_block3a56.port_b_first_address = 0;
defparam ram_block3a56.port_b_first_bit_number = 24;
defparam ram_block3a56.port_b_last_address = 8191;
defparam ram_block3a56.port_b_logical_ram_depth = 16384;
defparam ram_block3a56.port_b_logical_ram_width = 32;
defparam ram_block3a56.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_read_enable_clock = "clock1";
defparam ram_block3a56.port_b_write_enable_clock = "clock1";
defparam ram_block3a56.ram_block_type = "M9K";
defparam ram_block3a56.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y34_N0
cycloneive_ram_block ram_block3a24(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a24_PORTADATAOUT_bus),
	.portbdataout(ram_block3a24_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a24.clk0_core_clock_enable = "ena0";
defparam ram_block3a24.clk1_core_clock_enable = "ena1";
defparam ram_block3a24.data_interleave_offset_in_bits = 1;
defparam ram_block3a24.data_interleave_width_in_bits = 1;
defparam ram_block3a24.init_file = "meminit.hex";
defparam ram_block3a24.init_file_layout = "port_a";
defparam ram_block3a24.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a24.operation_mode = "bidir_dual_port";
defparam ram_block3a24.port_a_address_clear = "none";
defparam ram_block3a24.port_a_address_width = 13;
defparam ram_block3a24.port_a_byte_enable_clock = "none";
defparam ram_block3a24.port_a_data_out_clear = "none";
defparam ram_block3a24.port_a_data_out_clock = "none";
defparam ram_block3a24.port_a_data_width = 1;
defparam ram_block3a24.port_a_first_address = 0;
defparam ram_block3a24.port_a_first_bit_number = 24;
defparam ram_block3a24.port_a_last_address = 8191;
defparam ram_block3a24.port_a_logical_ram_depth = 16384;
defparam ram_block3a24.port_a_logical_ram_width = 32;
defparam ram_block3a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_address_clear = "none";
defparam ram_block3a24.port_b_address_clock = "clock1";
defparam ram_block3a24.port_b_address_width = 13;
defparam ram_block3a24.port_b_data_in_clock = "clock1";
defparam ram_block3a24.port_b_data_out_clear = "none";
defparam ram_block3a24.port_b_data_out_clock = "none";
defparam ram_block3a24.port_b_data_width = 1;
defparam ram_block3a24.port_b_first_address = 0;
defparam ram_block3a24.port_b_first_bit_number = 24;
defparam ram_block3a24.port_b_last_address = 8191;
defparam ram_block3a24.port_b_logical_ram_depth = 16384;
defparam ram_block3a24.port_b_logical_ram_width = 32;
defparam ram_block3a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_read_enable_clock = "clock1";
defparam ram_block3a24.port_b_write_enable_clock = "clock1";
defparam ram_block3a24.ram_block_type = "M9K";
defparam ram_block3a24.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000A000;
// synopsys translate_on

// Location: M9K_X64_Y46_N0
cycloneive_ram_block ram_block3a57(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a57_PORTADATAOUT_bus),
	.portbdataout(ram_block3a57_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a57.clk0_core_clock_enable = "ena0";
defparam ram_block3a57.clk1_core_clock_enable = "ena1";
defparam ram_block3a57.data_interleave_offset_in_bits = 1;
defparam ram_block3a57.data_interleave_width_in_bits = 1;
defparam ram_block3a57.init_file = "meminit.hex";
defparam ram_block3a57.init_file_layout = "port_a";
defparam ram_block3a57.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a57.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a57.operation_mode = "bidir_dual_port";
defparam ram_block3a57.port_a_address_clear = "none";
defparam ram_block3a57.port_a_address_width = 13;
defparam ram_block3a57.port_a_byte_enable_clock = "none";
defparam ram_block3a57.port_a_data_out_clear = "none";
defparam ram_block3a57.port_a_data_out_clock = "none";
defparam ram_block3a57.port_a_data_width = 1;
defparam ram_block3a57.port_a_first_address = 0;
defparam ram_block3a57.port_a_first_bit_number = 25;
defparam ram_block3a57.port_a_last_address = 8191;
defparam ram_block3a57.port_a_logical_ram_depth = 16384;
defparam ram_block3a57.port_a_logical_ram_width = 32;
defparam ram_block3a57.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_address_clear = "none";
defparam ram_block3a57.port_b_address_clock = "clock1";
defparam ram_block3a57.port_b_address_width = 13;
defparam ram_block3a57.port_b_data_in_clock = "clock1";
defparam ram_block3a57.port_b_data_out_clear = "none";
defparam ram_block3a57.port_b_data_out_clock = "none";
defparam ram_block3a57.port_b_data_width = 1;
defparam ram_block3a57.port_b_first_address = 0;
defparam ram_block3a57.port_b_first_bit_number = 25;
defparam ram_block3a57.port_b_last_address = 8191;
defparam ram_block3a57.port_b_logical_ram_depth = 16384;
defparam ram_block3a57.port_b_logical_ram_width = 32;
defparam ram_block3a57.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_read_enable_clock = "clock1";
defparam ram_block3a57.port_b_write_enable_clock = "clock1";
defparam ram_block3a57.ram_block_type = "M9K";
defparam ram_block3a57.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y42_N0
cycloneive_ram_block ram_block3a25(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a25_PORTADATAOUT_bus),
	.portbdataout(ram_block3a25_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a25.clk0_core_clock_enable = "ena0";
defparam ram_block3a25.clk1_core_clock_enable = "ena1";
defparam ram_block3a25.data_interleave_offset_in_bits = 1;
defparam ram_block3a25.data_interleave_width_in_bits = 1;
defparam ram_block3a25.init_file = "meminit.hex";
defparam ram_block3a25.init_file_layout = "port_a";
defparam ram_block3a25.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a25.operation_mode = "bidir_dual_port";
defparam ram_block3a25.port_a_address_clear = "none";
defparam ram_block3a25.port_a_address_width = 13;
defparam ram_block3a25.port_a_byte_enable_clock = "none";
defparam ram_block3a25.port_a_data_out_clear = "none";
defparam ram_block3a25.port_a_data_out_clock = "none";
defparam ram_block3a25.port_a_data_width = 1;
defparam ram_block3a25.port_a_first_address = 0;
defparam ram_block3a25.port_a_first_bit_number = 25;
defparam ram_block3a25.port_a_last_address = 8191;
defparam ram_block3a25.port_a_logical_ram_depth = 16384;
defparam ram_block3a25.port_a_logical_ram_width = 32;
defparam ram_block3a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_address_clear = "none";
defparam ram_block3a25.port_b_address_clock = "clock1";
defparam ram_block3a25.port_b_address_width = 13;
defparam ram_block3a25.port_b_data_in_clock = "clock1";
defparam ram_block3a25.port_b_data_out_clear = "none";
defparam ram_block3a25.port_b_data_out_clock = "none";
defparam ram_block3a25.port_b_data_width = 1;
defparam ram_block3a25.port_b_first_address = 0;
defparam ram_block3a25.port_b_first_bit_number = 25;
defparam ram_block3a25.port_b_last_address = 8191;
defparam ram_block3a25.port_b_logical_ram_depth = 16384;
defparam ram_block3a25.port_b_logical_ram_width = 32;
defparam ram_block3a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_read_enable_clock = "clock1";
defparam ram_block3a25.port_b_write_enable_clock = "clock1";
defparam ram_block3a25.ram_block_type = "M9K";
defparam ram_block3a25.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFE0000;
// synopsys translate_on

// Location: M9K_X51_Y40_N0
cycloneive_ram_block ram_block3a58(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a58_PORTADATAOUT_bus),
	.portbdataout(ram_block3a58_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a58.clk0_core_clock_enable = "ena0";
defparam ram_block3a58.clk1_core_clock_enable = "ena1";
defparam ram_block3a58.data_interleave_offset_in_bits = 1;
defparam ram_block3a58.data_interleave_width_in_bits = 1;
defparam ram_block3a58.init_file = "meminit.hex";
defparam ram_block3a58.init_file_layout = "port_a";
defparam ram_block3a58.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a58.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a58.operation_mode = "bidir_dual_port";
defparam ram_block3a58.port_a_address_clear = "none";
defparam ram_block3a58.port_a_address_width = 13;
defparam ram_block3a58.port_a_byte_enable_clock = "none";
defparam ram_block3a58.port_a_data_out_clear = "none";
defparam ram_block3a58.port_a_data_out_clock = "none";
defparam ram_block3a58.port_a_data_width = 1;
defparam ram_block3a58.port_a_first_address = 0;
defparam ram_block3a58.port_a_first_bit_number = 26;
defparam ram_block3a58.port_a_last_address = 8191;
defparam ram_block3a58.port_a_logical_ram_depth = 16384;
defparam ram_block3a58.port_a_logical_ram_width = 32;
defparam ram_block3a58.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_address_clear = "none";
defparam ram_block3a58.port_b_address_clock = "clock1";
defparam ram_block3a58.port_b_address_width = 13;
defparam ram_block3a58.port_b_data_in_clock = "clock1";
defparam ram_block3a58.port_b_data_out_clear = "none";
defparam ram_block3a58.port_b_data_out_clock = "none";
defparam ram_block3a58.port_b_data_width = 1;
defparam ram_block3a58.port_b_first_address = 0;
defparam ram_block3a58.port_b_first_bit_number = 26;
defparam ram_block3a58.port_b_last_address = 8191;
defparam ram_block3a58.port_b_logical_ram_depth = 16384;
defparam ram_block3a58.port_b_logical_ram_width = 32;
defparam ram_block3a58.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_read_enable_clock = "clock1";
defparam ram_block3a58.port_b_write_enable_clock = "clock1";
defparam ram_block3a58.ram_block_type = "M9K";
defparam ram_block3a58.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y44_N0
cycloneive_ram_block ram_block3a26(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a26_PORTADATAOUT_bus),
	.portbdataout(ram_block3a26_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a26.clk0_core_clock_enable = "ena0";
defparam ram_block3a26.clk1_core_clock_enable = "ena1";
defparam ram_block3a26.data_interleave_offset_in_bits = 1;
defparam ram_block3a26.data_interleave_width_in_bits = 1;
defparam ram_block3a26.init_file = "meminit.hex";
defparam ram_block3a26.init_file_layout = "port_a";
defparam ram_block3a26.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a26.operation_mode = "bidir_dual_port";
defparam ram_block3a26.port_a_address_clear = "none";
defparam ram_block3a26.port_a_address_width = 13;
defparam ram_block3a26.port_a_byte_enable_clock = "none";
defparam ram_block3a26.port_a_data_out_clear = "none";
defparam ram_block3a26.port_a_data_out_clock = "none";
defparam ram_block3a26.port_a_data_width = 1;
defparam ram_block3a26.port_a_first_address = 0;
defparam ram_block3a26.port_a_first_bit_number = 26;
defparam ram_block3a26.port_a_last_address = 8191;
defparam ram_block3a26.port_a_logical_ram_depth = 16384;
defparam ram_block3a26.port_a_logical_ram_width = 32;
defparam ram_block3a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_address_clear = "none";
defparam ram_block3a26.port_b_address_clock = "clock1";
defparam ram_block3a26.port_b_address_width = 13;
defparam ram_block3a26.port_b_data_in_clock = "clock1";
defparam ram_block3a26.port_b_data_out_clear = "none";
defparam ram_block3a26.port_b_data_out_clock = "none";
defparam ram_block3a26.port_b_data_width = 1;
defparam ram_block3a26.port_b_first_address = 0;
defparam ram_block3a26.port_b_first_bit_number = 26;
defparam ram_block3a26.port_b_last_address = 8191;
defparam ram_block3a26.port_b_logical_ram_depth = 16384;
defparam ram_block3a26.port_b_logical_ram_width = 32;
defparam ram_block3a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_read_enable_clock = "clock1";
defparam ram_block3a26.port_b_write_enable_clock = "clock1";
defparam ram_block3a26.ram_block_type = "M9K";
defparam ram_block3a26.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFE510F;
// synopsys translate_on

// Location: M9K_X51_Y46_N0
cycloneive_ram_block ram_block3a59(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a59_PORTADATAOUT_bus),
	.portbdataout(ram_block3a59_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a59.clk0_core_clock_enable = "ena0";
defparam ram_block3a59.clk1_core_clock_enable = "ena1";
defparam ram_block3a59.data_interleave_offset_in_bits = 1;
defparam ram_block3a59.data_interleave_width_in_bits = 1;
defparam ram_block3a59.init_file = "meminit.hex";
defparam ram_block3a59.init_file_layout = "port_a";
defparam ram_block3a59.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a59.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a59.operation_mode = "bidir_dual_port";
defparam ram_block3a59.port_a_address_clear = "none";
defparam ram_block3a59.port_a_address_width = 13;
defparam ram_block3a59.port_a_byte_enable_clock = "none";
defparam ram_block3a59.port_a_data_out_clear = "none";
defparam ram_block3a59.port_a_data_out_clock = "none";
defparam ram_block3a59.port_a_data_width = 1;
defparam ram_block3a59.port_a_first_address = 0;
defparam ram_block3a59.port_a_first_bit_number = 27;
defparam ram_block3a59.port_a_last_address = 8191;
defparam ram_block3a59.port_a_logical_ram_depth = 16384;
defparam ram_block3a59.port_a_logical_ram_width = 32;
defparam ram_block3a59.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_address_clear = "none";
defparam ram_block3a59.port_b_address_clock = "clock1";
defparam ram_block3a59.port_b_address_width = 13;
defparam ram_block3a59.port_b_data_in_clock = "clock1";
defparam ram_block3a59.port_b_data_out_clear = "none";
defparam ram_block3a59.port_b_data_out_clock = "none";
defparam ram_block3a59.port_b_data_width = 1;
defparam ram_block3a59.port_b_first_address = 0;
defparam ram_block3a59.port_b_first_bit_number = 27;
defparam ram_block3a59.port_b_last_address = 8191;
defparam ram_block3a59.port_b_logical_ram_depth = 16384;
defparam ram_block3a59.port_b_logical_ram_width = 32;
defparam ram_block3a59.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_read_enable_clock = "clock1";
defparam ram_block3a59.port_b_write_enable_clock = "clock1";
defparam ram_block3a59.ram_block_type = "M9K";
defparam ram_block3a59.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y43_N0
cycloneive_ram_block ram_block3a27(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a27_PORTADATAOUT_bus),
	.portbdataout(ram_block3a27_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a27.clk0_core_clock_enable = "ena0";
defparam ram_block3a27.clk1_core_clock_enable = "ena1";
defparam ram_block3a27.data_interleave_offset_in_bits = 1;
defparam ram_block3a27.data_interleave_width_in_bits = 1;
defparam ram_block3a27.init_file = "meminit.hex";
defparam ram_block3a27.init_file_layout = "port_a";
defparam ram_block3a27.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a27.operation_mode = "bidir_dual_port";
defparam ram_block3a27.port_a_address_clear = "none";
defparam ram_block3a27.port_a_address_width = 13;
defparam ram_block3a27.port_a_byte_enable_clock = "none";
defparam ram_block3a27.port_a_data_out_clear = "none";
defparam ram_block3a27.port_a_data_out_clock = "none";
defparam ram_block3a27.port_a_data_width = 1;
defparam ram_block3a27.port_a_first_address = 0;
defparam ram_block3a27.port_a_first_bit_number = 27;
defparam ram_block3a27.port_a_last_address = 8191;
defparam ram_block3a27.port_a_logical_ram_depth = 16384;
defparam ram_block3a27.port_a_logical_ram_width = 32;
defparam ram_block3a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_address_clear = "none";
defparam ram_block3a27.port_b_address_clock = "clock1";
defparam ram_block3a27.port_b_address_width = 13;
defparam ram_block3a27.port_b_data_in_clock = "clock1";
defparam ram_block3a27.port_b_data_out_clear = "none";
defparam ram_block3a27.port_b_data_out_clock = "none";
defparam ram_block3a27.port_b_data_width = 1;
defparam ram_block3a27.port_b_first_address = 0;
defparam ram_block3a27.port_b_first_bit_number = 27;
defparam ram_block3a27.port_b_last_address = 8191;
defparam ram_block3a27.port_b_logical_ram_depth = 16384;
defparam ram_block3a27.port_b_logical_ram_width = 32;
defparam ram_block3a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_read_enable_clock = "clock1";
defparam ram_block3a27.port_b_write_enable_clock = "clock1";
defparam ram_block3a27.ram_block_type = "M9K";
defparam ram_block3a27.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFE0800;
// synopsys translate_on

// Location: M9K_X64_Y40_N0
cycloneive_ram_block ram_block3a60(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a60_PORTADATAOUT_bus),
	.portbdataout(ram_block3a60_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a60.clk0_core_clock_enable = "ena0";
defparam ram_block3a60.clk1_core_clock_enable = "ena1";
defparam ram_block3a60.data_interleave_offset_in_bits = 1;
defparam ram_block3a60.data_interleave_width_in_bits = 1;
defparam ram_block3a60.init_file = "meminit.hex";
defparam ram_block3a60.init_file_layout = "port_a";
defparam ram_block3a60.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a60.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a60.operation_mode = "bidir_dual_port";
defparam ram_block3a60.port_a_address_clear = "none";
defparam ram_block3a60.port_a_address_width = 13;
defparam ram_block3a60.port_a_byte_enable_clock = "none";
defparam ram_block3a60.port_a_data_out_clear = "none";
defparam ram_block3a60.port_a_data_out_clock = "none";
defparam ram_block3a60.port_a_data_width = 1;
defparam ram_block3a60.port_a_first_address = 0;
defparam ram_block3a60.port_a_first_bit_number = 28;
defparam ram_block3a60.port_a_last_address = 8191;
defparam ram_block3a60.port_a_logical_ram_depth = 16384;
defparam ram_block3a60.port_a_logical_ram_width = 32;
defparam ram_block3a60.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_address_clear = "none";
defparam ram_block3a60.port_b_address_clock = "clock1";
defparam ram_block3a60.port_b_address_width = 13;
defparam ram_block3a60.port_b_data_in_clock = "clock1";
defparam ram_block3a60.port_b_data_out_clear = "none";
defparam ram_block3a60.port_b_data_out_clock = "none";
defparam ram_block3a60.port_b_data_width = 1;
defparam ram_block3a60.port_b_first_address = 0;
defparam ram_block3a60.port_b_first_bit_number = 28;
defparam ram_block3a60.port_b_last_address = 8191;
defparam ram_block3a60.port_b_logical_ram_depth = 16384;
defparam ram_block3a60.port_b_logical_ram_width = 32;
defparam ram_block3a60.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_read_enable_clock = "clock1";
defparam ram_block3a60.port_b_write_enable_clock = "clock1";
defparam ram_block3a60.ram_block_type = "M9K";
defparam ram_block3a60.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y47_N0
cycloneive_ram_block ram_block3a28(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a28_PORTADATAOUT_bus),
	.portbdataout(ram_block3a28_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a28.clk0_core_clock_enable = "ena0";
defparam ram_block3a28.clk1_core_clock_enable = "ena1";
defparam ram_block3a28.data_interleave_offset_in_bits = 1;
defparam ram_block3a28.data_interleave_width_in_bits = 1;
defparam ram_block3a28.init_file = "meminit.hex";
defparam ram_block3a28.init_file_layout = "port_a";
defparam ram_block3a28.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a28.operation_mode = "bidir_dual_port";
defparam ram_block3a28.port_a_address_clear = "none";
defparam ram_block3a28.port_a_address_width = 13;
defparam ram_block3a28.port_a_byte_enable_clock = "none";
defparam ram_block3a28.port_a_data_out_clear = "none";
defparam ram_block3a28.port_a_data_out_clock = "none";
defparam ram_block3a28.port_a_data_width = 1;
defparam ram_block3a28.port_a_first_address = 0;
defparam ram_block3a28.port_a_first_bit_number = 28;
defparam ram_block3a28.port_a_last_address = 8191;
defparam ram_block3a28.port_a_logical_ram_depth = 16384;
defparam ram_block3a28.port_a_logical_ram_width = 32;
defparam ram_block3a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_address_clear = "none";
defparam ram_block3a28.port_b_address_clock = "clock1";
defparam ram_block3a28.port_b_address_width = 13;
defparam ram_block3a28.port_b_data_in_clock = "clock1";
defparam ram_block3a28.port_b_data_out_clear = "none";
defparam ram_block3a28.port_b_data_out_clock = "none";
defparam ram_block3a28.port_b_data_width = 1;
defparam ram_block3a28.port_b_first_address = 0;
defparam ram_block3a28.port_b_first_bit_number = 28;
defparam ram_block3a28.port_b_last_address = 8191;
defparam ram_block3a28.port_b_logical_ram_depth = 16384;
defparam ram_block3a28.port_b_logical_ram_width = 32;
defparam ram_block3a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_read_enable_clock = "clock1";
defparam ram_block3a28.port_b_write_enable_clock = "clock1";
defparam ram_block3a28.ram_block_type = "M9K";
defparam ram_block3a28.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000584F;
// synopsys translate_on

// Location: M9K_X64_Y30_N0
cycloneive_ram_block ram_block3a61(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a61_PORTADATAOUT_bus),
	.portbdataout(ram_block3a61_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a61.clk0_core_clock_enable = "ena0";
defparam ram_block3a61.clk1_core_clock_enable = "ena1";
defparam ram_block3a61.data_interleave_offset_in_bits = 1;
defparam ram_block3a61.data_interleave_width_in_bits = 1;
defparam ram_block3a61.init_file = "meminit.hex";
defparam ram_block3a61.init_file_layout = "port_a";
defparam ram_block3a61.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a61.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a61.operation_mode = "bidir_dual_port";
defparam ram_block3a61.port_a_address_clear = "none";
defparam ram_block3a61.port_a_address_width = 13;
defparam ram_block3a61.port_a_byte_enable_clock = "none";
defparam ram_block3a61.port_a_data_out_clear = "none";
defparam ram_block3a61.port_a_data_out_clock = "none";
defparam ram_block3a61.port_a_data_width = 1;
defparam ram_block3a61.port_a_first_address = 0;
defparam ram_block3a61.port_a_first_bit_number = 29;
defparam ram_block3a61.port_a_last_address = 8191;
defparam ram_block3a61.port_a_logical_ram_depth = 16384;
defparam ram_block3a61.port_a_logical_ram_width = 32;
defparam ram_block3a61.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_address_clear = "none";
defparam ram_block3a61.port_b_address_clock = "clock1";
defparam ram_block3a61.port_b_address_width = 13;
defparam ram_block3a61.port_b_data_in_clock = "clock1";
defparam ram_block3a61.port_b_data_out_clear = "none";
defparam ram_block3a61.port_b_data_out_clock = "none";
defparam ram_block3a61.port_b_data_width = 1;
defparam ram_block3a61.port_b_first_address = 0;
defparam ram_block3a61.port_b_first_bit_number = 29;
defparam ram_block3a61.port_b_last_address = 8191;
defparam ram_block3a61.port_b_logical_ram_depth = 16384;
defparam ram_block3a61.port_b_logical_ram_width = 32;
defparam ram_block3a61.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_read_enable_clock = "clock1";
defparam ram_block3a61.port_b_write_enable_clock = "clock1";
defparam ram_block3a61.ram_block_type = "M9K";
defparam ram_block3a61.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y25_N0
cycloneive_ram_block ram_block3a29(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a29_PORTADATAOUT_bus),
	.portbdataout(ram_block3a29_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a29.clk0_core_clock_enable = "ena0";
defparam ram_block3a29.clk1_core_clock_enable = "ena1";
defparam ram_block3a29.data_interleave_offset_in_bits = 1;
defparam ram_block3a29.data_interleave_width_in_bits = 1;
defparam ram_block3a29.init_file = "meminit.hex";
defparam ram_block3a29.init_file_layout = "port_a";
defparam ram_block3a29.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a29.operation_mode = "bidir_dual_port";
defparam ram_block3a29.port_a_address_clear = "none";
defparam ram_block3a29.port_a_address_width = 13;
defparam ram_block3a29.port_a_byte_enable_clock = "none";
defparam ram_block3a29.port_a_data_out_clear = "none";
defparam ram_block3a29.port_a_data_out_clock = "none";
defparam ram_block3a29.port_a_data_width = 1;
defparam ram_block3a29.port_a_first_address = 0;
defparam ram_block3a29.port_a_first_bit_number = 29;
defparam ram_block3a29.port_a_last_address = 8191;
defparam ram_block3a29.port_a_logical_ram_depth = 16384;
defparam ram_block3a29.port_a_logical_ram_width = 32;
defparam ram_block3a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_address_clear = "none";
defparam ram_block3a29.port_b_address_clock = "clock1";
defparam ram_block3a29.port_b_address_width = 13;
defparam ram_block3a29.port_b_data_in_clock = "clock1";
defparam ram_block3a29.port_b_data_out_clear = "none";
defparam ram_block3a29.port_b_data_out_clock = "none";
defparam ram_block3a29.port_b_data_width = 1;
defparam ram_block3a29.port_b_first_address = 0;
defparam ram_block3a29.port_b_first_bit_number = 29;
defparam ram_block3a29.port_b_last_address = 8191;
defparam ram_block3a29.port_b_logical_ram_depth = 16384;
defparam ram_block3a29.port_b_logical_ram_width = 32;
defparam ram_block3a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_read_enable_clock = "clock1";
defparam ram_block3a29.port_b_write_enable_clock = "clock1";
defparam ram_block3a29.ram_block_type = "M9K";
defparam ram_block3a29.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFE594F;
// synopsys translate_on

// Location: M9K_X64_Y38_N0
cycloneive_ram_block ram_block3a62(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a62_PORTADATAOUT_bus),
	.portbdataout(ram_block3a62_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a62.clk0_core_clock_enable = "ena0";
defparam ram_block3a62.clk1_core_clock_enable = "ena1";
defparam ram_block3a62.data_interleave_offset_in_bits = 1;
defparam ram_block3a62.data_interleave_width_in_bits = 1;
defparam ram_block3a62.init_file = "meminit.hex";
defparam ram_block3a62.init_file_layout = "port_a";
defparam ram_block3a62.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a62.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a62.operation_mode = "bidir_dual_port";
defparam ram_block3a62.port_a_address_clear = "none";
defparam ram_block3a62.port_a_address_width = 13;
defparam ram_block3a62.port_a_byte_enable_clock = "none";
defparam ram_block3a62.port_a_data_out_clear = "none";
defparam ram_block3a62.port_a_data_out_clock = "none";
defparam ram_block3a62.port_a_data_width = 1;
defparam ram_block3a62.port_a_first_address = 0;
defparam ram_block3a62.port_a_first_bit_number = 30;
defparam ram_block3a62.port_a_last_address = 8191;
defparam ram_block3a62.port_a_logical_ram_depth = 16384;
defparam ram_block3a62.port_a_logical_ram_width = 32;
defparam ram_block3a62.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_address_clear = "none";
defparam ram_block3a62.port_b_address_clock = "clock1";
defparam ram_block3a62.port_b_address_width = 13;
defparam ram_block3a62.port_b_data_in_clock = "clock1";
defparam ram_block3a62.port_b_data_out_clear = "none";
defparam ram_block3a62.port_b_data_out_clock = "none";
defparam ram_block3a62.port_b_data_width = 1;
defparam ram_block3a62.port_b_first_address = 0;
defparam ram_block3a62.port_b_first_bit_number = 30;
defparam ram_block3a62.port_b_last_address = 8191;
defparam ram_block3a62.port_b_logical_ram_depth = 16384;
defparam ram_block3a62.port_b_logical_ram_width = 32;
defparam ram_block3a62.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_read_enable_clock = "clock1";
defparam ram_block3a62.port_b_write_enable_clock = "clock1";
defparam ram_block3a62.ram_block_type = "M9K";
defparam ram_block3a62.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y27_N0
cycloneive_ram_block ram_block3a30(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a30_PORTADATAOUT_bus),
	.portbdataout(ram_block3a30_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a30.clk0_core_clock_enable = "ena0";
defparam ram_block3a30.clk1_core_clock_enable = "ena1";
defparam ram_block3a30.data_interleave_offset_in_bits = 1;
defparam ram_block3a30.data_interleave_width_in_bits = 1;
defparam ram_block3a30.init_file = "meminit.hex";
defparam ram_block3a30.init_file_layout = "port_a";
defparam ram_block3a30.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a30.operation_mode = "bidir_dual_port";
defparam ram_block3a30.port_a_address_clear = "none";
defparam ram_block3a30.port_a_address_width = 13;
defparam ram_block3a30.port_a_byte_enable_clock = "none";
defparam ram_block3a30.port_a_data_out_clear = "none";
defparam ram_block3a30.port_a_data_out_clock = "none";
defparam ram_block3a30.port_a_data_width = 1;
defparam ram_block3a30.port_a_first_address = 0;
defparam ram_block3a30.port_a_first_bit_number = 30;
defparam ram_block3a30.port_a_last_address = 8191;
defparam ram_block3a30.port_a_logical_ram_depth = 16384;
defparam ram_block3a30.port_a_logical_ram_width = 32;
defparam ram_block3a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_address_clear = "none";
defparam ram_block3a30.port_b_address_clock = "clock1";
defparam ram_block3a30.port_b_address_width = 13;
defparam ram_block3a30.port_b_data_in_clock = "clock1";
defparam ram_block3a30.port_b_data_out_clear = "none";
defparam ram_block3a30.port_b_data_out_clock = "none";
defparam ram_block3a30.port_b_data_width = 1;
defparam ram_block3a30.port_b_first_address = 0;
defparam ram_block3a30.port_b_first_bit_number = 30;
defparam ram_block3a30.port_b_last_address = 8191;
defparam ram_block3a30.port_b_logical_ram_depth = 16384;
defparam ram_block3a30.port_b_logical_ram_width = 32;
defparam ram_block3a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_read_enable_clock = "clock1";
defparam ram_block3a30.port_b_write_enable_clock = "clock1";
defparam ram_block3a30.ram_block_type = "M9K";
defparam ram_block3a30.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000;
// synopsys translate_on

// Location: M9K_X51_Y26_N0
cycloneive_ram_block ram_block3a63(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a63_PORTADATAOUT_bus),
	.portbdataout(ram_block3a63_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a63.clk0_core_clock_enable = "ena0";
defparam ram_block3a63.clk1_core_clock_enable = "ena1";
defparam ram_block3a63.data_interleave_offset_in_bits = 1;
defparam ram_block3a63.data_interleave_width_in_bits = 1;
defparam ram_block3a63.init_file = "meminit.hex";
defparam ram_block3a63.init_file_layout = "port_a";
defparam ram_block3a63.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a63.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a63.operation_mode = "bidir_dual_port";
defparam ram_block3a63.port_a_address_clear = "none";
defparam ram_block3a63.port_a_address_width = 13;
defparam ram_block3a63.port_a_byte_enable_clock = "none";
defparam ram_block3a63.port_a_data_out_clear = "none";
defparam ram_block3a63.port_a_data_out_clock = "none";
defparam ram_block3a63.port_a_data_width = 1;
defparam ram_block3a63.port_a_first_address = 0;
defparam ram_block3a63.port_a_first_bit_number = 31;
defparam ram_block3a63.port_a_last_address = 8191;
defparam ram_block3a63.port_a_logical_ram_depth = 16384;
defparam ram_block3a63.port_a_logical_ram_width = 32;
defparam ram_block3a63.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_address_clear = "none";
defparam ram_block3a63.port_b_address_clock = "clock1";
defparam ram_block3a63.port_b_address_width = 13;
defparam ram_block3a63.port_b_data_in_clock = "clock1";
defparam ram_block3a63.port_b_data_out_clear = "none";
defparam ram_block3a63.port_b_data_out_clock = "none";
defparam ram_block3a63.port_b_data_width = 1;
defparam ram_block3a63.port_b_first_address = 0;
defparam ram_block3a63.port_b_first_bit_number = 31;
defparam ram_block3a63.port_b_last_address = 8191;
defparam ram_block3a63.port_b_logical_ram_depth = 16384;
defparam ram_block3a63.port_b_logical_ram_width = 32;
defparam ram_block3a63.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_read_enable_clock = "clock1";
defparam ram_block3a63.port_b_write_enable_clock = "clock1";
defparam ram_block3a63.ram_block_type = "M9K";
defparam ram_block3a63.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y26_N0
cycloneive_ram_block ram_block3a31(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a31_PORTADATAOUT_bus),
	.portbdataout(ram_block3a31_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a31.clk0_core_clock_enable = "ena0";
defparam ram_block3a31.clk1_core_clock_enable = "ena1";
defparam ram_block3a31.data_interleave_offset_in_bits = 1;
defparam ram_block3a31.data_interleave_width_in_bits = 1;
defparam ram_block3a31.init_file = "meminit.hex";
defparam ram_block3a31.init_file_layout = "port_a";
defparam ram_block3a31.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a31.operation_mode = "bidir_dual_port";
defparam ram_block3a31.port_a_address_clear = "none";
defparam ram_block3a31.port_a_address_width = 13;
defparam ram_block3a31.port_a_byte_enable_clock = "none";
defparam ram_block3a31.port_a_data_out_clear = "none";
defparam ram_block3a31.port_a_data_out_clock = "none";
defparam ram_block3a31.port_a_data_width = 1;
defparam ram_block3a31.port_a_first_address = 0;
defparam ram_block3a31.port_a_first_bit_number = 31;
defparam ram_block3a31.port_a_last_address = 8191;
defparam ram_block3a31.port_a_logical_ram_depth = 16384;
defparam ram_block3a31.port_a_logical_ram_width = 32;
defparam ram_block3a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_address_clear = "none";
defparam ram_block3a31.port_b_address_clock = "clock1";
defparam ram_block3a31.port_b_address_width = 13;
defparam ram_block3a31.port_b_data_in_clock = "clock1";
defparam ram_block3a31.port_b_data_out_clear = "none";
defparam ram_block3a31.port_b_data_out_clock = "none";
defparam ram_block3a31.port_b_data_width = 1;
defparam ram_block3a31.port_b_first_address = 0;
defparam ram_block3a31.port_b_first_bit_number = 31;
defparam ram_block3a31.port_b_last_address = 8191;
defparam ram_block3a31.port_b_logical_ram_depth = 16384;
defparam ram_block3a31.port_b_logical_ram_width = 32;
defparam ram_block3a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_read_enable_clock = "clock1";
defparam ram_block3a31.port_b_write_enable_clock = "clock1";
defparam ram_block3a31.ram_block_type = "M9K";
defparam ram_block3a31.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFE0000;
// synopsys translate_on

// Location: FF_X59_Y34_N5
dffeas \address_reg_a[0] (
	.clk(clock0),
	.d(gnd),
	.asdata(ramaddr1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_a_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_a[0] .is_wysiwyg = "true";
defparam \address_reg_a[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N7
dffeas \address_reg_b[0] (
	.clk(clock1),
	.d(\address_reg_b[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_b_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_b[0] .is_wysiwyg = "true";
defparam \address_reg_b[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N6
cycloneive_lcell_comb \address_reg_b[0]~feeder (
// Equation(s):
// \address_reg_b[0]~feeder_combout  = ram_rom_addr_reg_13

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_13),
	.cin(gnd),
	.combout(\address_reg_b[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \address_reg_b[0]~feeder .lut_mask = 16'hFF00;
defparam \address_reg_b[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa (
	ramaddr,
	ramWEN,
	always1,
	eq_node_1,
	eq_node_0,
	devpor,
	devclrn,
	devoe);
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	eq_node_1;
output 	eq_node_0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X65_Y34_N4
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (!\ramWEN~0_combout  & (always1 & !\ramaddr~29_combout ))

	.dataa(gnd),
	.datab(ramWEN),
	.datac(always1),
	.datad(ramaddr),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h0030;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N30
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (!\ramWEN~0_combout  & (always1 & \ramaddr~29_combout ))

	.dataa(gnd),
	.datab(ramWEN),
	.datac(always1),
	.datad(ramaddr),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h3000;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa_1 (
	ram_rom_addr_reg_13,
	sdr,
	eq_node_1,
	eq_node_0,
	irf_reg_2_1,
	state_5,
	devpor,
	devclrn,
	devoe);
input 	ram_rom_addr_reg_13;
input 	sdr;
output 	eq_node_1;
output 	eq_node_0;
input 	irf_reg_2_1;
input 	state_5;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X42_Y41_N28
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (sdr & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & (ram_rom_addr_reg_13 & \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q )))

	.dataa(sdr),
	.datab(state_5),
	.datac(ram_rom_addr_reg_13),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h8000;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N22
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (sdr & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & (!ram_rom_addr_reg_13 & \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q )))

	.dataa(sdr),
	.datab(state_5),
	.datac(ram_rom_addr_reg_13),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h0800;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_mod_ram_rom (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg1,
	ram_rom_data_reg_0,
	ram_rom_addr_reg_13,
	ram_rom_addr_reg_0,
	ram_rom_addr_reg_1,
	ram_rom_addr_reg_2,
	ram_rom_addr_reg_3,
	ram_rom_addr_reg_4,
	ram_rom_addr_reg_5,
	ram_rom_addr_reg_6,
	ram_rom_addr_reg_7,
	ram_rom_addr_reg_8,
	ram_rom_addr_reg_9,
	ram_rom_addr_reg_10,
	ram_rom_addr_reg_11,
	ram_rom_addr_reg_12,
	ram_rom_data_reg_1,
	ram_rom_data_reg_2,
	ram_rom_data_reg_3,
	ram_rom_data_reg_4,
	ram_rom_data_reg_5,
	ram_rom_data_reg_6,
	ram_rom_data_reg_7,
	ram_rom_data_reg_8,
	ram_rom_data_reg_9,
	ram_rom_data_reg_10,
	ram_rom_data_reg_11,
	ram_rom_data_reg_12,
	ram_rom_data_reg_13,
	ram_rom_data_reg_14,
	ram_rom_data_reg_15,
	ram_rom_data_reg_16,
	ram_rom_data_reg_17,
	ram_rom_data_reg_18,
	ram_rom_data_reg_19,
	ram_rom_data_reg_20,
	ram_rom_data_reg_21,
	ram_rom_data_reg_22,
	ram_rom_data_reg_23,
	ram_rom_data_reg_24,
	ram_rom_data_reg_25,
	ram_rom_data_reg_26,
	ram_rom_data_reg_27,
	ram_rom_data_reg_28,
	ram_rom_data_reg_29,
	ram_rom_data_reg_30,
	ram_rom_data_reg_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	sdr,
	address_reg_b_0,
	altera_internal_jtag,
	state_4,
	ir_in,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_4_1,
	node_ena_1,
	clr,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	raw_tck,
	devpor,
	devclrn,
	devoe);
input 	ram_block3a32;
input 	ram_block3a0;
input 	ram_block3a33;
input 	ram_block3a1;
input 	ram_block3a34;
input 	ram_block3a2;
input 	ram_block3a35;
input 	ram_block3a3;
input 	ram_block3a36;
input 	ram_block3a4;
input 	ram_block3a37;
input 	ram_block3a5;
input 	ram_block3a38;
input 	ram_block3a6;
input 	ram_block3a39;
input 	ram_block3a7;
input 	ram_block3a40;
input 	ram_block3a8;
input 	ram_block3a41;
input 	ram_block3a9;
input 	ram_block3a42;
input 	ram_block3a10;
input 	ram_block3a43;
input 	ram_block3a11;
input 	ram_block3a44;
input 	ram_block3a12;
input 	ram_block3a45;
input 	ram_block3a13;
input 	ram_block3a46;
input 	ram_block3a14;
input 	ram_block3a47;
input 	ram_block3a15;
input 	ram_block3a48;
input 	ram_block3a16;
input 	ram_block3a49;
input 	ram_block3a17;
input 	ram_block3a50;
input 	ram_block3a18;
input 	ram_block3a51;
input 	ram_block3a19;
input 	ram_block3a52;
input 	ram_block3a20;
input 	ram_block3a53;
input 	ram_block3a21;
input 	ram_block3a54;
input 	ram_block3a22;
input 	ram_block3a55;
input 	ram_block3a23;
input 	ram_block3a56;
input 	ram_block3a24;
input 	ram_block3a57;
input 	ram_block3a25;
input 	ram_block3a58;
input 	ram_block3a26;
input 	ram_block3a59;
input 	ram_block3a27;
input 	ram_block3a60;
input 	ram_block3a28;
input 	ram_block3a61;
input 	ram_block3a29;
input 	ram_block3a62;
input 	ram_block3a30;
input 	ram_block3a63;
input 	ram_block3a31;
output 	is_in_use_reg1;
output 	ram_rom_data_reg_0;
output 	ram_rom_addr_reg_13;
output 	ram_rom_addr_reg_0;
output 	ram_rom_addr_reg_1;
output 	ram_rom_addr_reg_2;
output 	ram_rom_addr_reg_3;
output 	ram_rom_addr_reg_4;
output 	ram_rom_addr_reg_5;
output 	ram_rom_addr_reg_6;
output 	ram_rom_addr_reg_7;
output 	ram_rom_addr_reg_8;
output 	ram_rom_addr_reg_9;
output 	ram_rom_addr_reg_10;
output 	ram_rom_addr_reg_11;
output 	ram_rom_addr_reg_12;
output 	ram_rom_data_reg_1;
output 	ram_rom_data_reg_2;
output 	ram_rom_data_reg_3;
output 	ram_rom_data_reg_4;
output 	ram_rom_data_reg_5;
output 	ram_rom_data_reg_6;
output 	ram_rom_data_reg_7;
output 	ram_rom_data_reg_8;
output 	ram_rom_data_reg_9;
output 	ram_rom_data_reg_10;
output 	ram_rom_data_reg_11;
output 	ram_rom_data_reg_12;
output 	ram_rom_data_reg_13;
output 	ram_rom_data_reg_14;
output 	ram_rom_data_reg_15;
output 	ram_rom_data_reg_16;
output 	ram_rom_data_reg_17;
output 	ram_rom_data_reg_18;
output 	ram_rom_data_reg_19;
output 	ram_rom_data_reg_20;
output 	ram_rom_data_reg_21;
output 	ram_rom_data_reg_22;
output 	ram_rom_data_reg_23;
output 	ram_rom_data_reg_24;
output 	ram_rom_data_reg_25;
output 	ram_rom_data_reg_26;
output 	ram_rom_data_reg_27;
output 	ram_rom_data_reg_28;
output 	ram_rom_data_reg_29;
output 	ram_rom_data_reg_30;
output 	ram_rom_data_reg_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
output 	sdr;
input 	address_reg_b_0;
input 	altera_internal_jtag;
input 	state_4;
input 	[4:0] ir_in;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	raw_tck;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~2_combout ;
wire \Add1~6_combout ;
wire \ram_rom_data_shift_cntr_reg[3]~8_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~12_combout ;
wire \is_in_use_reg~0_combout ;
wire \ram_rom_data_reg[0]~0_combout ;
wire \Add1~0_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~4_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~11_combout ;
wire \ram_rom_data_shift_cntr_reg[0]~6_combout ;
wire \Add1~1 ;
wire \Add1~3 ;
wire \Add1~4_combout ;
wire \ram_rom_data_shift_cntr_reg[2]~9_combout ;
wire \Add1~5 ;
wire \Add1~7 ;
wire \Add1~8_combout ;
wire \ram_rom_data_shift_cntr_reg[4]~7_combout ;
wire \Add1~9 ;
wire \Add1~10_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~10_combout ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \ram_rom_data_shift_cntr_reg[1]~5_combout ;
wire \process_0~2_combout ;
wire \ram_rom_data_reg[0]~32_combout ;
wire \ram_rom_addr_reg[0]~15 ;
wire \ram_rom_addr_reg[1]~17 ;
wire \ram_rom_addr_reg[2]~19 ;
wire \ram_rom_addr_reg[3]~21 ;
wire \ram_rom_addr_reg[4]~23 ;
wire \ram_rom_addr_reg[5]~25 ;
wire \ram_rom_addr_reg[6]~27 ;
wire \ram_rom_addr_reg[7]~29 ;
wire \ram_rom_addr_reg[8]~31 ;
wire \ram_rom_addr_reg[9]~33 ;
wire \ram_rom_addr_reg[10]~35 ;
wire \ram_rom_addr_reg[11]~37 ;
wire \ram_rom_addr_reg[12]~39 ;
wire \ram_rom_addr_reg[13]~40_combout ;
wire \process_0~3_combout ;
wire \ram_rom_addr_reg[5]~42_combout ;
wire \ram_rom_addr_reg[5]~43_combout ;
wire \ram_rom_addr_reg[0]~14_combout ;
wire \ram_rom_addr_reg[1]~16_combout ;
wire \ram_rom_addr_reg[2]~18_combout ;
wire \ram_rom_addr_reg[3]~20_combout ;
wire \ram_rom_addr_reg[4]~22_combout ;
wire \ram_rom_addr_reg[5]~24_combout ;
wire \ram_rom_addr_reg[6]~26_combout ;
wire \ram_rom_addr_reg[7]~28_combout ;
wire \ram_rom_addr_reg[8]~30_combout ;
wire \ram_rom_addr_reg[9]~32_combout ;
wire \ram_rom_addr_reg[10]~34_combout ;
wire \ram_rom_addr_reg[11]~36_combout ;
wire \ram_rom_addr_reg[12]~38_combout ;
wire \ram_rom_data_reg[1]~1_combout ;
wire \ram_rom_data_reg[2]~2_combout ;
wire \ram_rom_data_reg[3]~3_combout ;
wire \ram_rom_data_reg[4]~4_combout ;
wire \ram_rom_data_reg[5]~5_combout ;
wire \ram_rom_data_reg[6]~6_combout ;
wire \ram_rom_data_reg[7]~7_combout ;
wire \ram_rom_data_reg[8]~8_combout ;
wire \ram_rom_data_reg[9]~9_combout ;
wire \ram_rom_data_reg[10]~10_combout ;
wire \ram_rom_data_reg[11]~11_combout ;
wire \ram_rom_data_reg[12]~12_combout ;
wire \ram_rom_data_reg[13]~13_combout ;
wire \ram_rom_data_reg[14]~14_combout ;
wire \ram_rom_data_reg[15]~15_combout ;
wire \ram_rom_data_reg[16]~16_combout ;
wire \ram_rom_data_reg[17]~17_combout ;
wire \ram_rom_data_reg[18]~18_combout ;
wire \ram_rom_data_reg[19]~19_combout ;
wire \ram_rom_data_reg[20]~20_combout ;
wire \ram_rom_data_reg[21]~21_combout ;
wire \ram_rom_data_reg[22]~22_combout ;
wire \ram_rom_data_reg[23]~23_combout ;
wire \ram_rom_data_reg[24]~24_combout ;
wire \ram_rom_data_reg[25]~25_combout ;
wire \ram_rom_data_reg[26]~26_combout ;
wire \ram_rom_data_reg[27]~27_combout ;
wire \ram_rom_data_reg[28]~28_combout ;
wire \ram_rom_data_reg[29]~29_combout ;
wire \ram_rom_data_reg[30]~30_combout ;
wire \ram_rom_data_reg[31]~31_combout ;
wire \ir_loaded_address_reg[0]~feeder_combout ;
wire \process_0~0_combout ;
wire \process_0~1_combout ;
wire \ir_loaded_address_reg[1]~feeder_combout ;
wire \ir_loaded_address_reg[3]~feeder_combout ;
wire \bypass_reg_out~0_combout ;
wire \bypass_reg_out~q ;
wire \tdo~0_combout ;
wire [5:0] ram_rom_data_shift_cntr_reg;
wire [3:0] \ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR ;


sld_rom_sr \ram_rom_logic_gen:name_gen:info_rom_sr (
	.WORD_SR_0(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.sdr(sdr),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.TCK(raw_tck),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X41_Y42_N14
cycloneive_lcell_comb \Add1~2 (
	.dataa(ram_rom_data_shift_cntr_reg[1]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h5A5F;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X41_Y42_N18
cycloneive_lcell_comb \Add1~6 (
	.dataa(ram_rom_data_shift_cntr_reg[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h5A5F;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X41_Y42_N31
dffeas \ram_rom_data_shift_cntr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[3]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y42_N30
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[3]~8 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~6_combout ),
	.datac(ram_rom_data_shift_cntr_reg[3]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3]~8 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[3]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y42_N6
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~12 (
	.dataa(ram_rom_data_shift_cntr_reg[1]),
	.datab(\Equal1~0_combout ),
	.datac(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datad(ram_rom_data_shift_cntr_reg[0]),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~12 .lut_mask = 16'h8F0F;
defparam \ram_rom_data_shift_cntr_reg[5]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y41_N25
dffeas is_in_use_reg(
	.clk(raw_tck),
	.d(\is_in_use_reg~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(ir_in[0]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(is_in_use_reg1),
	.prn(vcc));
// synopsys translate_off
defparam is_in_use_reg.is_wysiwyg = "true";
defparam is_in_use_reg.power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N21
dffeas \ram_rom_data_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[0]~0_combout ),
	.asdata(ram_rom_data_reg_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N31
dffeas \ram_rom_addr_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[13]~40_combout ),
	.asdata(altera_internal_jtag),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N5
dffeas \ram_rom_addr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[0]~14_combout ),
	.asdata(ram_rom_addr_reg_1),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N7
dffeas \ram_rom_addr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[1]~16_combout ),
	.asdata(ram_rom_addr_reg_2),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N9
dffeas \ram_rom_addr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[2]~18_combout ),
	.asdata(ram_rom_addr_reg_3),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N11
dffeas \ram_rom_addr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[3]~20_combout ),
	.asdata(ram_rom_addr_reg_4),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N13
dffeas \ram_rom_addr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[4]~22_combout ),
	.asdata(ram_rom_addr_reg_5),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N15
dffeas \ram_rom_addr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[5]~24_combout ),
	.asdata(ram_rom_addr_reg_6),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N17
dffeas \ram_rom_addr_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[6]~26_combout ),
	.asdata(ram_rom_addr_reg_7),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N19
dffeas \ram_rom_addr_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[7]~28_combout ),
	.asdata(ram_rom_addr_reg_8),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N21
dffeas \ram_rom_addr_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[8]~30_combout ),
	.asdata(ram_rom_addr_reg_9),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N23
dffeas \ram_rom_addr_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[9]~32_combout ),
	.asdata(ram_rom_addr_reg_10),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N25
dffeas \ram_rom_addr_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[10]~34_combout ),
	.asdata(ram_rom_addr_reg_11),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N27
dffeas \ram_rom_addr_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[11]~36_combout ),
	.asdata(ram_rom_addr_reg_12),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N29
dffeas \ram_rom_addr_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[12]~38_combout ),
	.asdata(ram_rom_addr_reg_13),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N27
dffeas \ram_rom_data_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[1]~1_combout ),
	.asdata(ram_rom_data_reg_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N13
dffeas \ram_rom_data_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[2]~2_combout ),
	.asdata(ram_rom_data_reg_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N11
dffeas \ram_rom_data_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[3]~3_combout ),
	.asdata(ram_rom_data_reg_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N9
dffeas \ram_rom_data_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[4]~4_combout ),
	.asdata(ram_rom_data_reg_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N13
dffeas \ram_rom_data_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[5]~5_combout ),
	.asdata(ram_rom_data_reg_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N31
dffeas \ram_rom_data_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[6]~6_combout ),
	.asdata(ram_rom_data_reg_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N17
dffeas \ram_rom_data_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[7]~7_combout ),
	.asdata(ram_rom_data_reg_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N7
dffeas \ram_rom_data_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[8]~8_combout ),
	.asdata(ram_rom_data_reg_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N5
dffeas \ram_rom_data_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[9]~9_combout ),
	.asdata(ram_rom_data_reg_10),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N17
dffeas \ram_rom_data_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[10]~10_combout ),
	.asdata(ram_rom_data_reg_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N23
dffeas \ram_rom_data_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[11]~11_combout ),
	.asdata(ram_rom_data_reg_12),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N27
dffeas \ram_rom_data_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[12]~12_combout ),
	.asdata(ram_rom_data_reg_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N9
dffeas \ram_rom_data_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[13]~13_combout ),
	.asdata(ram_rom_data_reg_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N21
dffeas \ram_rom_data_reg[14] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[14]~14_combout ),
	.asdata(ram_rom_data_reg_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_14),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[14] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N11
dffeas \ram_rom_data_reg[15] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[15]~15_combout ),
	.asdata(ram_rom_data_reg_16),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_15),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[15] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N29
dffeas \ram_rom_data_reg[16] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[16]~16_combout ),
	.asdata(ram_rom_data_reg_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_16),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[16] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N31
dffeas \ram_rom_data_reg[17] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[17]~17_combout ),
	.asdata(ram_rom_data_reg_18),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_17),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[17] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N25
dffeas \ram_rom_data_reg[18] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[18]~18_combout ),
	.asdata(ram_rom_data_reg_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_18),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[18] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N15
dffeas \ram_rom_data_reg[19] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[19]~19_combout ),
	.asdata(ram_rom_data_reg_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_19),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[19] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N13
dffeas \ram_rom_data_reg[20] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[20]~20_combout ),
	.asdata(ram_rom_data_reg_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_20),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[20] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N15
dffeas \ram_rom_data_reg[21] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[21]~21_combout ),
	.asdata(ram_rom_data_reg_22),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_21),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[21] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N29
dffeas \ram_rom_data_reg[22] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[22]~22_combout ),
	.asdata(ram_rom_data_reg_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_22),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[22] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N31
dffeas \ram_rom_data_reg[23] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[23]~23_combout ),
	.asdata(ram_rom_data_reg_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_23),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[23] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y39_N15
dffeas \ram_rom_data_reg[24] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[24]~24_combout ),
	.asdata(ram_rom_data_reg_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_24),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[24] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N21
dffeas \ram_rom_data_reg[25] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[25]~25_combout ),
	.asdata(ram_rom_data_reg_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_25),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[25] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N11
dffeas \ram_rom_data_reg[26] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[26]~26_combout ),
	.asdata(ram_rom_data_reg_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_26),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[26] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N9
dffeas \ram_rom_data_reg[27] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[27]~27_combout ),
	.asdata(ram_rom_data_reg_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_27),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[27] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N23
dffeas \ram_rom_data_reg[28] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[28]~28_combout ),
	.asdata(ram_rom_data_reg_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_28),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[28] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N5
dffeas \ram_rom_data_reg[29] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[29]~29_combout ),
	.asdata(ram_rom_data_reg_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_29),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[29] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N19
dffeas \ram_rom_data_reg[30] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[30]~30_combout ),
	.asdata(ram_rom_data_reg_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_30),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[30] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N25
dffeas \ram_rom_data_reg[31] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[31]~31_combout ),
	.asdata(altera_internal_jtag),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_31),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[31] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y42_N21
dffeas \ir_loaded_address_reg[0] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[0] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y41_N15
dffeas \ir_loaded_address_reg[1] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[1] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y42_N31
dffeas \ir_loaded_address_reg[2] (
	.clk(raw_tck),
	.d(gnd),
	.asdata(ram_rom_addr_reg_2),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[2] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y42_N5
dffeas \ir_loaded_address_reg[3] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[3] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N4
cycloneive_lcell_comb \tdo~1 (
	.dataa(gnd),
	.datab(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.datac(ir_in[0]),
	.datad(\tdo~0_combout ),
	.cin(gnd),
	.combout(tdo),
	.cout());
// synopsys translate_off
defparam \tdo~1 .lut_mask = 16'hCFC0;
defparam \tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N6
cycloneive_lcell_comb \sdr~0 (
	.dataa(gnd),
	.datab(node_ena_1),
	.datac(virtual_ir_scan_reg),
	.datad(gnd),
	.cin(gnd),
	.combout(sdr),
	.cout());
// synopsys translate_off
defparam \sdr~0 .lut_mask = 16'h0C0C;
defparam \sdr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N24
cycloneive_lcell_comb \is_in_use_reg~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(is_in_use_reg1),
	.datad(irf_reg_4_1),
	.cin(gnd),
	.combout(\is_in_use_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \is_in_use_reg~0 .lut_mask = 16'h00F0;
defparam \is_in_use_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N20
cycloneive_lcell_comb \ram_rom_data_reg[0]~0 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a32),
	.datac(gnd),
	.datad(ram_block3a0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[0]~0 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y42_N12
cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h33CC;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N30
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~4 (
	.dataa(irf_reg_1_1),
	.datab(sdr),
	.datac(state_4),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~4 .lut_mask = 16'hC080;
defparam \ram_rom_data_shift_cntr_reg[5]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y42_N28
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~11 (
	.dataa(ram_rom_data_shift_cntr_reg[1]),
	.datab(\Equal1~0_combout ),
	.datac(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datad(ram_rom_data_shift_cntr_reg[0]),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~11 .lut_mask = 16'h070F;
defparam \ram_rom_data_shift_cntr_reg[5]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y42_N2
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[0]~6 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~0_combout ),
	.datac(ram_rom_data_shift_cntr_reg[0]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0]~6 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[0]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y42_N3
dffeas \ram_rom_data_shift_cntr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[0]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y42_N16
cycloneive_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'hC30C;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X41_Y42_N0
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[2]~9 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~4_combout ),
	.datac(ram_rom_data_shift_cntr_reg[2]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2]~9 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[2]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y42_N1
dffeas \ram_rom_data_shift_cntr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[2]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y42_N20
cycloneive_lcell_comb \Add1~8 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'hC30C;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X41_Y42_N4
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[4]~7 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~8_combout ),
	.datac(ram_rom_data_shift_cntr_reg[4]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4]~7 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[4]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y42_N5
dffeas \ram_rom_data_shift_cntr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[4]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y42_N22
cycloneive_lcell_comb \Add1~10 (
	.dataa(ram_rom_data_shift_cntr_reg[5]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h5A5A;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X41_Y42_N26
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~10 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~10_combout ),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~10 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[5]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y42_N27
dffeas \ram_rom_data_shift_cntr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[5]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y42_N24
cycloneive_lcell_comb \Equal1~0 (
	.dataa(ram_rom_data_shift_cntr_reg[3]),
	.datab(ram_rom_data_shift_cntr_reg[4]),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(ram_rom_data_shift_cntr_reg[2]),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h0800;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y42_N10
cycloneive_lcell_comb \Equal1~1 (
	.dataa(gnd),
	.datab(\Equal1~0_combout ),
	.datac(gnd),
	.datad(ram_rom_data_shift_cntr_reg[0]),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~1 .lut_mask = 16'hCC00;
defparam \Equal1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y42_N8
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[1]~5 (
	.dataa(\Add1~2_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1]~5 .lut_mask = 16'h08B8;
defparam \ram_rom_data_shift_cntr_reg[1]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y42_N9
dffeas \ram_rom_data_shift_cntr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[1]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N12
cycloneive_lcell_comb \process_0~2 (
	.dataa(\Equal1~1_combout ),
	.datab(ram_rom_data_shift_cntr_reg[1]),
	.datac(ir_in[3]),
	.datad(irf_reg_1_1),
	.cin(gnd),
	.combout(\process_0~2_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~2 .lut_mask = 16'h070F;
defparam \process_0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N24
cycloneive_lcell_comb \ram_rom_data_reg[0]~32 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\process_0~2_combout ),
	.datad(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_reg[0]~32_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[0]~32 .lut_mask = 16'hFF0F;
defparam \ram_rom_data_reg[0]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N4
cycloneive_lcell_comb \ram_rom_addr_reg[0]~14 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[0]~14_combout ),
	.cout(\ram_rom_addr_reg[0]~15 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[0]~14 .lut_mask = 16'h33CC;
defparam \ram_rom_addr_reg[0]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N6
cycloneive_lcell_comb \ram_rom_addr_reg[1]~16 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[0]~15 ),
	.combout(\ram_rom_addr_reg[1]~16_combout ),
	.cout(\ram_rom_addr_reg[1]~17 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[1]~16 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[1]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N8
cycloneive_lcell_comb \ram_rom_addr_reg[2]~18 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[1]~17 ),
	.combout(\ram_rom_addr_reg[2]~18_combout ),
	.cout(\ram_rom_addr_reg[2]~19 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[2]~18 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[2]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N10
cycloneive_lcell_comb \ram_rom_addr_reg[3]~20 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[2]~19 ),
	.combout(\ram_rom_addr_reg[3]~20_combout ),
	.cout(\ram_rom_addr_reg[3]~21 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[3]~20 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[3]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N12
cycloneive_lcell_comb \ram_rom_addr_reg[4]~22 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[3]~21 ),
	.combout(\ram_rom_addr_reg[4]~22_combout ),
	.cout(\ram_rom_addr_reg[4]~23 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[4]~22 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[4]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N14
cycloneive_lcell_comb \ram_rom_addr_reg[5]~24 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[4]~23 ),
	.combout(\ram_rom_addr_reg[5]~24_combout ),
	.cout(\ram_rom_addr_reg[5]~25 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[5]~24 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[5]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N16
cycloneive_lcell_comb \ram_rom_addr_reg[6]~26 (
	.dataa(ram_rom_addr_reg_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[5]~25 ),
	.combout(\ram_rom_addr_reg[6]~26_combout ),
	.cout(\ram_rom_addr_reg[6]~27 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[6]~26 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[6]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N18
cycloneive_lcell_comb \ram_rom_addr_reg[7]~28 (
	.dataa(ram_rom_addr_reg_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[6]~27 ),
	.combout(\ram_rom_addr_reg[7]~28_combout ),
	.cout(\ram_rom_addr_reg[7]~29 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[7]~28 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[7]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N20
cycloneive_lcell_comb \ram_rom_addr_reg[8]~30 (
	.dataa(ram_rom_addr_reg_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[7]~29 ),
	.combout(\ram_rom_addr_reg[8]~30_combout ),
	.cout(\ram_rom_addr_reg[8]~31 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[8]~30 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[8]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N22
cycloneive_lcell_comb \ram_rom_addr_reg[9]~32 (
	.dataa(ram_rom_addr_reg_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[8]~31 ),
	.combout(\ram_rom_addr_reg[9]~32_combout ),
	.cout(\ram_rom_addr_reg[9]~33 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[9]~32 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[9]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N24
cycloneive_lcell_comb \ram_rom_addr_reg[10]~34 (
	.dataa(ram_rom_addr_reg_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[9]~33 ),
	.combout(\ram_rom_addr_reg[10]~34_combout ),
	.cout(\ram_rom_addr_reg[10]~35 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[10]~34 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[10]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N26
cycloneive_lcell_comb \ram_rom_addr_reg[11]~36 (
	.dataa(ram_rom_addr_reg_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[10]~35 ),
	.combout(\ram_rom_addr_reg[11]~36_combout ),
	.cout(\ram_rom_addr_reg[11]~37 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[11]~36 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[11]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N28
cycloneive_lcell_comb \ram_rom_addr_reg[12]~38 (
	.dataa(ram_rom_addr_reg_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[11]~37 ),
	.combout(\ram_rom_addr_reg[12]~38_combout ),
	.cout(\ram_rom_addr_reg[12]~39 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[12]~38 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[12]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N30
cycloneive_lcell_comb \ram_rom_addr_reg[13]~40 (
	.dataa(ram_rom_addr_reg_13),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\ram_rom_addr_reg[12]~39 ),
	.combout(\ram_rom_addr_reg[13]~40_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[13]~40 .lut_mask = 16'h5A5A;
defparam \ram_rom_addr_reg[13]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N8
cycloneive_lcell_comb \process_0~3 (
	.dataa(state_4),
	.datab(ir_in[3]),
	.datac(node_ena_1),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\process_0~3_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~3 .lut_mask = 16'h0080;
defparam \process_0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N2
cycloneive_lcell_comb \ram_rom_addr_reg[5]~42 (
	.dataa(irf_reg_1_1),
	.datab(\process_0~3_combout ),
	.datac(\Equal1~1_combout ),
	.datad(ram_rom_data_shift_cntr_reg[1]),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[5]~42_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[5]~42 .lut_mask = 16'hCCEC;
defparam \ram_rom_addr_reg[5]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N16
cycloneive_lcell_comb \ram_rom_addr_reg[5]~43 (
	.dataa(sdr),
	.datab(\ram_rom_addr_reg[5]~42_combout ),
	.datac(state_8),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[5]~43_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[5]~43 .lut_mask = 16'hECCC;
defparam \ram_rom_addr_reg[5]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N26
cycloneive_lcell_comb \ram_rom_data_reg[1]~1 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a33),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_rom_data_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[1]~1 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N12
cycloneive_lcell_comb \ram_rom_data_reg[2]~2 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a2),
	.datac(gnd),
	.datad(ram_block3a34),
	.cin(gnd),
	.combout(\ram_rom_data_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[2]~2 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N10
cycloneive_lcell_comb \ram_rom_data_reg[3]~3 (
	.dataa(ram_block3a35),
	.datab(ram_block3a3),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[3]~3 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N8
cycloneive_lcell_comb \ram_rom_data_reg[4]~4 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a36),
	.datac(gnd),
	.datad(ram_block3a4),
	.cin(gnd),
	.combout(\ram_rom_data_reg[4]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[4]~4 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N12
cycloneive_lcell_comb \ram_rom_data_reg[5]~5 (
	.dataa(ram_block3a5),
	.datab(ram_block3a37),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[5]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[5]~5 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[5]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N30
cycloneive_lcell_comb \ram_rom_data_reg[6]~6 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a38),
	.datac(gnd),
	.datad(ram_block3a6),
	.cin(gnd),
	.combout(\ram_rom_data_reg[6]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[6]~6 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[6]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N16
cycloneive_lcell_comb \ram_rom_data_reg[7]~7 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a39),
	.datac(gnd),
	.datad(ram_block3a7),
	.cin(gnd),
	.combout(\ram_rom_data_reg[7]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[7]~7 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[7]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N6
cycloneive_lcell_comb \ram_rom_data_reg[8]~8 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a8),
	.datac(gnd),
	.datad(ram_block3a40),
	.cin(gnd),
	.combout(\ram_rom_data_reg[8]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[8]~8 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[8]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N4
cycloneive_lcell_comb \ram_rom_data_reg[9]~9 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a9),
	.datac(gnd),
	.datad(ram_block3a41),
	.cin(gnd),
	.combout(\ram_rom_data_reg[9]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[9]~9 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[9]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N16
cycloneive_lcell_comb \ram_rom_data_reg[10]~10 (
	.dataa(ram_block3a42),
	.datab(ram_block3a10),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[10]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[10]~10 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[10]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N22
cycloneive_lcell_comb \ram_rom_data_reg[11]~11 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a43),
	.datac(gnd),
	.datad(ram_block3a11),
	.cin(gnd),
	.combout(\ram_rom_data_reg[11]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[11]~11 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[11]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N26
cycloneive_lcell_comb \ram_rom_data_reg[12]~12 (
	.dataa(ram_block3a12),
	.datab(ram_block3a44),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[12]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[12]~12 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N8
cycloneive_lcell_comb \ram_rom_data_reg[13]~13 (
	.dataa(ram_block3a45),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a13),
	.cin(gnd),
	.combout(\ram_rom_data_reg[13]~13_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[13]~13 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[13]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N20
cycloneive_lcell_comb \ram_rom_data_reg[14]~14 (
	.dataa(ram_block3a46),
	.datab(ram_block3a14),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[14]~14_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[14]~14 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[14]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N10
cycloneive_lcell_comb \ram_rom_data_reg[15]~15 (
	.dataa(ram_block3a15),
	.datab(ram_block3a47),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[15]~15_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[15]~15 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[15]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N28
cycloneive_lcell_comb \ram_rom_data_reg[16]~16 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a16),
	.datac(gnd),
	.datad(ram_block3a48),
	.cin(gnd),
	.combout(\ram_rom_data_reg[16]~16_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[16]~16 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[16]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N30
cycloneive_lcell_comb \ram_rom_data_reg[17]~17 (
	.dataa(ram_block3a49),
	.datab(ram_block3a17),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[17]~17_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[17]~17 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[17]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N24
cycloneive_lcell_comb \ram_rom_data_reg[18]~18 (
	.dataa(ram_block3a18),
	.datab(ram_block3a50),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[18]~18_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[18]~18 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[18]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N14
cycloneive_lcell_comb \ram_rom_data_reg[19]~19 (
	.dataa(ram_block3a51),
	.datab(ram_block3a19),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[19]~19_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[19]~19 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[19]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N12
cycloneive_lcell_comb \ram_rom_data_reg[20]~20 (
	.dataa(ram_block3a20),
	.datab(ram_block3a52),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[20]~20_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[20]~20 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[20]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N14
cycloneive_lcell_comb \ram_rom_data_reg[21]~21 (
	.dataa(ram_block3a21),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a53),
	.cin(gnd),
	.combout(\ram_rom_data_reg[21]~21_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[21]~21 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[21]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N28
cycloneive_lcell_comb \ram_rom_data_reg[22]~22 (
	.dataa(ram_block3a54),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a22),
	.cin(gnd),
	.combout(\ram_rom_data_reg[22]~22_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[22]~22 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[22]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N30
cycloneive_lcell_comb \ram_rom_data_reg[23]~23 (
	.dataa(ram_block3a23),
	.datab(ram_block3a55),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[23]~23_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[23]~23 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[23]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y39_N14
cycloneive_lcell_comb \ram_rom_data_reg[24]~24 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a24),
	.datac(gnd),
	.datad(ram_block3a56),
	.cin(gnd),
	.combout(\ram_rom_data_reg[24]~24_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[24]~24 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[24]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N20
cycloneive_lcell_comb \ram_rom_data_reg[25]~25 (
	.dataa(ram_block3a25),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a57),
	.cin(gnd),
	.combout(\ram_rom_data_reg[25]~25_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[25]~25 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[25]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N10
cycloneive_lcell_comb \ram_rom_data_reg[26]~26 (
	.dataa(ram_block3a58),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a26),
	.cin(gnd),
	.combout(\ram_rom_data_reg[26]~26_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[26]~26 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[26]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N8
cycloneive_lcell_comb \ram_rom_data_reg[27]~27 (
	.dataa(ram_block3a59),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a27),
	.cin(gnd),
	.combout(\ram_rom_data_reg[27]~27_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[27]~27 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[27]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N22
cycloneive_lcell_comb \ram_rom_data_reg[28]~28 (
	.dataa(ram_block3a60),
	.datab(ram_block3a28),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[28]~28_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[28]~28 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[28]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N4
cycloneive_lcell_comb \ram_rom_data_reg[29]~29 (
	.dataa(ram_block3a29),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a61),
	.cin(gnd),
	.combout(\ram_rom_data_reg[29]~29_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[29]~29 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N18
cycloneive_lcell_comb \ram_rom_data_reg[30]~30 (
	.dataa(ram_block3a62),
	.datab(ram_block3a30),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[30]~30_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[30]~30 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N24
cycloneive_lcell_comb \ram_rom_data_reg[31]~31 (
	.dataa(ram_block3a31),
	.datab(ram_block3a63),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[31]~31_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[31]~31 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[31]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y42_N20
cycloneive_lcell_comb \ir_loaded_address_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_0),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N0
cycloneive_lcell_comb \process_0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ir_in[0]),
	.datad(irf_reg_4_1),
	.cin(gnd),
	.combout(\process_0~0_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~0 .lut_mask = 16'hFFF0;
defparam \process_0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N10
cycloneive_lcell_comb \process_0~1 (
	.dataa(virtual_ir_scan_reg),
	.datab(node_ena_1),
	.datac(ir_in[3]),
	.datad(state_5),
	.cin(gnd),
	.combout(\process_0~1_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~1 .lut_mask = 16'h4000;
defparam \process_0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N14
cycloneive_lcell_comb \ir_loaded_address_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_1),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y42_N4
cycloneive_lcell_comb \ir_loaded_address_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_3),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N20
cycloneive_lcell_comb \bypass_reg_out~0 (
	.dataa(gnd),
	.datab(node_ena_1),
	.datac(\bypass_reg_out~q ),
	.datad(altera_internal_jtag),
	.cin(gnd),
	.combout(\bypass_reg_out~0_combout ),
	.cout());
// synopsys translate_off
defparam \bypass_reg_out~0 .lut_mask = 16'hFC30;
defparam \bypass_reg_out~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y41_N21
dffeas bypass_reg_out(
	.clk(raw_tck),
	.d(\bypass_reg_out~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\bypass_reg_out~q ),
	.prn(vcc));
// synopsys translate_off
defparam bypass_reg_out.is_wysiwyg = "true";
defparam bypass_reg_out.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N18
cycloneive_lcell_comb \tdo~0 (
	.dataa(irf_reg_1_1),
	.datab(\bypass_reg_out~q ),
	.datac(ram_rom_data_reg_0),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(\tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \tdo~0 .lut_mask = 16'hF0E4;
defparam \tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_rom_sr (
	WORD_SR_0,
	sdr,
	altera_internal_jtag,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	TCK,
	devpor,
	devclrn,
	devoe);
output 	WORD_SR_0;
input 	sdr;
input 	altera_internal_jtag;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	TCK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \WORD_SR~3_combout ;
wire \word_counter[2]~13_combout ;
wire \WORD_SR~13_combout ;
wire \WORD_SR~14_combout ;
wire \WORD_SR~15_combout ;
wire \word_counter[0]~7_combout ;
wire \word_counter[2]~19_combout ;
wire \clear_signal~combout ;
wire \word_counter[2]~14_combout ;
wire \word_counter[0]~8 ;
wire \word_counter[1]~9_combout ;
wire \word_counter[1]~10 ;
wire \word_counter[2]~11_combout ;
wire \word_counter[2]~12 ;
wire \word_counter[3]~15_combout ;
wire \WORD_SR~2_combout ;
wire \WORD_SR~4_combout ;
wire \WORD_SR~10_combout ;
wire \WORD_SR~11_combout ;
wire \WORD_SR~12_combout ;
wire \WORD_SR[0]~6_combout ;
wire \word_counter[3]~16 ;
wire \word_counter[4]~17_combout ;
wire \WORD_SR~7_combout ;
wire \WORD_SR~8_combout ;
wire \WORD_SR~9_combout ;
wire \WORD_SR~5_combout ;
wire [4:0] word_counter;
wire [3:0] WORD_SR;


// Location: LCCOMB_X40_Y41_N10
cycloneive_lcell_comb \WORD_SR~3 (
	.dataa(word_counter[4]),
	.datab(word_counter[2]),
	.datac(word_counter[0]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~3_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~3 .lut_mask = 16'hAE02;
defparam \WORD_SR~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y41_N10
cycloneive_lcell_comb \word_counter[2]~13 (
	.dataa(word_counter[1]),
	.datab(word_counter[3]),
	.datac(word_counter[2]),
	.datad(word_counter[4]),
	.cin(gnd),
	.combout(\word_counter[2]~13_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[2]~13 .lut_mask = 16'hEFFF;
defparam \word_counter[2]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y41_N23
dffeas \WORD_SR[3] (
	.clk(TCK),
	.d(\WORD_SR~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[0]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[3]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[3] .is_wysiwyg = "true";
defparam \WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y41_N8
cycloneive_lcell_comb \WORD_SR~13 (
	.dataa(word_counter[1]),
	.datab(word_counter[3]),
	.datac(word_counter[2]),
	.datad(word_counter[4]),
	.cin(gnd),
	.combout(\WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~13 .lut_mask = 16'h0080;
defparam \WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y41_N18
cycloneive_lcell_comb \WORD_SR~14 (
	.dataa(altera_internal_jtag),
	.datab(state_4),
	.datac(\WORD_SR~13_combout ),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~14 .lut_mask = 16'h88B8;
defparam \WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y41_N22
cycloneive_lcell_comb \WORD_SR~15 (
	.dataa(state_8),
	.datab(gnd),
	.datac(virtual_ir_scan_reg),
	.datad(\WORD_SR~14_combout ),
	.cin(gnd),
	.combout(\WORD_SR~15_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~15 .lut_mask = 16'h5F00;
defparam \WORD_SR~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y41_N25
dffeas \WORD_SR[0] (
	.clk(TCK),
	.d(\WORD_SR~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[0]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR_0),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[0] .is_wysiwyg = "true";
defparam \WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y41_N22
cycloneive_lcell_comb \word_counter[0]~7 (
	.dataa(word_counter[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\word_counter[0]~7_combout ),
	.cout(\word_counter[0]~8 ));
// synopsys translate_off
defparam \word_counter[0]~7 .lut_mask = 16'h55AA;
defparam \word_counter[0]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y41_N20
cycloneive_lcell_comb \word_counter[2]~19 (
	.dataa(\word_counter[2]~13_combout ),
	.datab(word_counter[0]),
	.datac(virtual_ir_scan_reg),
	.datad(state_8),
	.cin(gnd),
	.combout(\word_counter[2]~19_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[2]~19 .lut_mask = 16'hF111;
defparam \word_counter[2]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y41_N0
cycloneive_lcell_comb clear_signal(
	.dataa(gnd),
	.datab(gnd),
	.datac(virtual_ir_scan_reg),
	.datad(state_8),
	.cin(gnd),
	.combout(\clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam clear_signal.lut_mask = 16'hF000;
defparam clear_signal.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y41_N12
cycloneive_lcell_comb \word_counter[2]~14 (
	.dataa(sdr),
	.datab(state_4),
	.datac(state_3),
	.datad(\clear_signal~combout ),
	.cin(gnd),
	.combout(\word_counter[2]~14_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[2]~14 .lut_mask = 16'hFF20;
defparam \word_counter[2]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y41_N23
dffeas \word_counter[0] (
	.clk(TCK),
	.d(\word_counter[0]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[2]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[2]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[0]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[0] .is_wysiwyg = "true";
defparam \word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y41_N24
cycloneive_lcell_comb \word_counter[1]~9 (
	.dataa(gnd),
	.datab(word_counter[1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[0]~8 ),
	.combout(\word_counter[1]~9_combout ),
	.cout(\word_counter[1]~10 ));
// synopsys translate_off
defparam \word_counter[1]~9 .lut_mask = 16'h3C3F;
defparam \word_counter[1]~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X40_Y41_N25
dffeas \word_counter[1] (
	.clk(TCK),
	.d(\word_counter[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[2]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[2]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[1]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[1] .is_wysiwyg = "true";
defparam \word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y41_N26
cycloneive_lcell_comb \word_counter[2]~11 (
	.dataa(gnd),
	.datab(word_counter[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[1]~10 ),
	.combout(\word_counter[2]~11_combout ),
	.cout(\word_counter[2]~12 ));
// synopsys translate_off
defparam \word_counter[2]~11 .lut_mask = 16'hC30C;
defparam \word_counter[2]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X40_Y41_N27
dffeas \word_counter[2] (
	.clk(TCK),
	.d(\word_counter[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[2]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[2]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[2]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[2] .is_wysiwyg = "true";
defparam \word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y41_N28
cycloneive_lcell_comb \word_counter[3]~15 (
	.dataa(gnd),
	.datab(word_counter[3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[2]~12 ),
	.combout(\word_counter[3]~15_combout ),
	.cout(\word_counter[3]~16 ));
// synopsys translate_off
defparam \word_counter[3]~15 .lut_mask = 16'h3C3F;
defparam \word_counter[3]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X40_Y41_N29
dffeas \word_counter[3] (
	.clk(TCK),
	.d(\word_counter[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[2]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[2]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[3]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[3] .is_wysiwyg = "true";
defparam \word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y41_N12
cycloneive_lcell_comb \WORD_SR~2 (
	.dataa(word_counter[4]),
	.datab(word_counter[1]),
	.datac(word_counter[2]),
	.datad(word_counter[3]),
	.cin(gnd),
	.combout(\WORD_SR~2_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~2 .lut_mask = 16'h5003;
defparam \WORD_SR~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y41_N16
cycloneive_lcell_comb \WORD_SR~4 (
	.dataa(\WORD_SR~3_combout ),
	.datab(gnd),
	.datac(word_counter[0]),
	.datad(\WORD_SR~2_combout ),
	.cin(gnd),
	.combout(\WORD_SR~4_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~4 .lut_mask = 16'hAAA0;
defparam \WORD_SR~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y41_N2
cycloneive_lcell_comb \WORD_SR~10 (
	.dataa(word_counter[4]),
	.datab(word_counter[2]),
	.datac(word_counter[0]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~10 .lut_mask = 16'hE2AE;
defparam \WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y41_N0
cycloneive_lcell_comb \WORD_SR~11 (
	.dataa(gnd),
	.datab(\WORD_SR~10_combout ),
	.datac(word_counter[0]),
	.datad(\WORD_SR~2_combout ),
	.cin(gnd),
	.combout(\WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~11 .lut_mask = 16'hC3C0;
defparam \WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y41_N28
cycloneive_lcell_comb \WORD_SR~12 (
	.dataa(WORD_SR[3]),
	.datab(state_4),
	.datac(\WORD_SR~11_combout ),
	.datad(\clear_signal~combout ),
	.cin(gnd),
	.combout(\WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~12 .lut_mask = 16'h00B8;
defparam \WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y41_N26
cycloneive_lcell_comb \WORD_SR[0]~6 (
	.dataa(sdr),
	.datab(state_4),
	.datac(state_3),
	.datad(\clear_signal~combout ),
	.cin(gnd),
	.combout(\WORD_SR[0]~6_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR[0]~6 .lut_mask = 16'hFFA8;
defparam \WORD_SR[0]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y41_N29
dffeas \WORD_SR[2] (
	.clk(TCK),
	.d(\WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[0]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[2]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[2] .is_wysiwyg = "true";
defparam \WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y41_N30
cycloneive_lcell_comb \word_counter[4]~17 (
	.dataa(word_counter[4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\word_counter[3]~16 ),
	.combout(\word_counter[4]~17_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[4]~17 .lut_mask = 16'hA5A5;
defparam \word_counter[4]~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X40_Y41_N31
dffeas \word_counter[4] (
	.clk(TCK),
	.d(\word_counter[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[2]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[2]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[4]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[4] .is_wysiwyg = "true";
defparam \word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y41_N16
cycloneive_lcell_comb \WORD_SR~7 (
	.dataa(word_counter[1]),
	.datab(word_counter[4]),
	.datac(state_4),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~7 .lut_mask = 16'h000B;
defparam \WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y41_N30
cycloneive_lcell_comb \WORD_SR~8 (
	.dataa(gnd),
	.datab(word_counter[3]),
	.datac(word_counter[2]),
	.datad(\WORD_SR~7_combout ),
	.cin(gnd),
	.combout(\WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~8 .lut_mask = 16'h0300;
defparam \WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y41_N14
cycloneive_lcell_comb \WORD_SR~9 (
	.dataa(state_4),
	.datab(WORD_SR[2]),
	.datac(\WORD_SR~8_combout ),
	.datad(\clear_signal~combout ),
	.cin(gnd),
	.combout(\WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~9 .lut_mask = 16'h00F8;
defparam \WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y41_N15
dffeas \WORD_SR[1] (
	.clk(TCK),
	.d(\WORD_SR~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[0]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[1]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[1] .is_wysiwyg = "true";
defparam \WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y41_N24
cycloneive_lcell_comb \WORD_SR~5 (
	.dataa(\WORD_SR~4_combout ),
	.datab(state_4),
	.datac(WORD_SR[1]),
	.datad(\clear_signal~combout ),
	.cin(gnd),
	.combout(\WORD_SR~5_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~5 .lut_mask = 16'h00E2;
defparam \WORD_SR~5 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module singlecycle (
	PC_29,
	PC_28,
	PC_31,
	PC_30,
	dpifhalt,
	PC_1,
	daddr_1,
	reg_WEN,
	reg_REN,
	PC_0,
	daddr_0,
	daddr_3,
	PC_3,
	daddr_2,
	PC_2,
	daddr_5,
	PC_5,
	PC_4,
	daddr_4,
	PC_7,
	daddr_7,
	daddr_6,
	PC_6,
	daddr_9,
	PC_9,
	daddr_8,
	PC_8,
	daddr_11,
	PC_11,
	daddr_10,
	PC_10,
	PC_13,
	daddr_13,
	daddr_12,
	PC_12,
	daddr_15,
	PC_15,
	daddr_14,
	PC_14,
	daddr_17,
	PC_17,
	PC_16,
	daddr_16,
	daddr_19,
	PC_19,
	daddr_18,
	PC_18,
	PC_21,
	daddr_21,
	daddr_20,
	PC_20,
	daddr_23,
	PC_23,
	daddr_22,
	PC_22,
	daddr_25,
	PC_25,
	daddr_24,
	PC_24,
	PC_27,
	daddr_27,
	daddr_26,
	PC_26,
	daddr_29,
	daddr_28,
	daddr_31,
	daddr_30,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	Mux63,
	Mux631,
	dcifimemload_20,
	Mux32,
	Mux321,
	Mux33,
	Mux331,
	Mux34,
	Mux341,
	Mux35,
	Mux351,
	Mux36,
	Mux361,
	Mux37,
	Mux371,
	Mux38,
	Mux381,
	Mux39,
	Mux391,
	Mux40,
	Mux401,
	Mux41,
	Mux411,
	Mux42,
	Mux421,
	Mux43,
	Mux431,
	Mux44,
	Mux441,
	Mux45,
	Mux451,
	Mux46,
	Mux461,
	Mux47,
	Mux471,
	Mux48,
	Mux481,
	Mux49,
	Mux491,
	Mux50,
	Mux501,
	Mux51,
	Mux511,
	Mux52,
	Mux521,
	Mux53,
	Mux531,
	Mux54,
	Mux541,
	Mux55,
	Mux551,
	Mux56,
	Mux561,
	Mux57,
	Mux571,
	Mux58,
	Mux581,
	Mux59,
	Mux591,
	Mux60,
	Mux601,
	Mux61,
	Mux611,
	Mux62,
	Mux621,
	nRST,
	CLK,
	nRST1,
	devpor,
	devclrn,
	devoe);
output 	PC_29;
output 	PC_28;
output 	PC_31;
output 	PC_30;
output 	dpifhalt;
output 	PC_1;
output 	daddr_1;
output 	reg_WEN;
output 	reg_REN;
output 	PC_0;
output 	daddr_0;
output 	daddr_3;
output 	PC_3;
output 	daddr_2;
output 	PC_2;
output 	daddr_5;
output 	PC_5;
output 	PC_4;
output 	daddr_4;
output 	PC_7;
output 	daddr_7;
output 	daddr_6;
output 	PC_6;
output 	daddr_9;
output 	PC_9;
output 	daddr_8;
output 	PC_8;
output 	daddr_11;
output 	PC_11;
output 	daddr_10;
output 	PC_10;
output 	PC_13;
output 	daddr_13;
output 	daddr_12;
output 	PC_12;
output 	daddr_15;
output 	PC_15;
output 	daddr_14;
output 	PC_14;
output 	daddr_17;
output 	PC_17;
output 	PC_16;
output 	daddr_16;
output 	daddr_19;
output 	PC_19;
output 	daddr_18;
output 	PC_18;
output 	PC_21;
output 	daddr_21;
output 	daddr_20;
output 	PC_20;
output 	daddr_23;
output 	PC_23;
output 	daddr_22;
output 	PC_22;
output 	daddr_25;
output 	PC_25;
output 	daddr_24;
output 	PC_24;
output 	PC_27;
output 	daddr_27;
output 	daddr_26;
output 	PC_26;
output 	daddr_29;
output 	daddr_28;
output 	daddr_31;
output 	daddr_30;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
output 	Mux63;
output 	Mux631;
output 	dcifimemload_20;
output 	Mux32;
output 	Mux321;
output 	Mux33;
output 	Mux331;
output 	Mux34;
output 	Mux341;
output 	Mux35;
output 	Mux351;
output 	Mux36;
output 	Mux361;
output 	Mux37;
output 	Mux371;
output 	Mux38;
output 	Mux381;
output 	Mux39;
output 	Mux391;
output 	Mux40;
output 	Mux401;
output 	Mux41;
output 	Mux411;
output 	Mux42;
output 	Mux421;
output 	Mux43;
output 	Mux431;
output 	Mux44;
output 	Mux441;
output 	Mux45;
output 	Mux451;
output 	Mux46;
output 	Mux461;
output 	Mux47;
output 	Mux471;
output 	Mux48;
output 	Mux481;
output 	Mux49;
output 	Mux491;
output 	Mux50;
output 	Mux501;
output 	Mux51;
output 	Mux511;
output 	Mux52;
output 	Mux521;
output 	Mux53;
output 	Mux531;
output 	Mux54;
output 	Mux541;
output 	Mux55;
output 	Mux551;
output 	Mux56;
output 	Mux561;
output 	Mux57;
output 	Mux571;
output 	Mux58;
output 	Mux581;
output 	Mux59;
output 	Mux591;
output 	Mux60;
output 	Mux601;
output 	Mux61;
output 	Mux611;
output 	Mux62;
output 	Mux621;
input 	nRST;
input 	CLK;
input 	nRST1;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \CC|ccif.iwait[0]~0_combout ;
wire \CM|dcif.imemload[30]~0_combout ;
wire \CM|dcif.imemload[31]~1_combout ;
wire \CM|dcif.imemload[27]~2_combout ;
wire \CM|dcif.imemload[26]~3_combout ;
wire \CM|dcif.imemload[29]~4_combout ;
wire \CM|dcif.imemload[28]~5_combout ;
wire \CM|dcif.imemload[19]~6_combout ;
wire \CM|dcif.imemload[18]~7_combout ;
wire \CM|dcif.imemload[16]~8_combout ;
wire \CM|dcif.imemload[17]~9_combout ;
wire \CM|dcif.imemload[24]~11_combout ;
wire \CM|dcif.imemload[23]~12_combout ;
wire \CM|dcif.imemload[21]~13_combout ;
wire \CM|dcif.imemload[22]~14_combout ;
wire \CM|dcif.imemload[25]~15_combout ;
wire \CM|dcif.imemload[3]~16_combout ;
wire \CM|dcif.imemload[4]~17_combout ;
wire \CM|dcif.imemload[2]~18_combout ;
wire \CM|dcif.imemload[5]~19_combout ;
wire \CM|dcif.imemload[0]~20_combout ;
wire \CM|dcif.imemload[1]~21_combout ;
wire \CM|dcif.imemload[15]~22_combout ;
wire \CM|dcif.imemload[14]~23_combout ;
wire \CM|dcif.imemload[13]~24_combout ;
wire \CM|dcif.imemload[12]~25_combout ;
wire \CM|dcif.imemload[11]~26_combout ;
wire \CM|dcif.imemload[10]~27_combout ;
wire \CM|dcif.imemload[9]~28_combout ;
wire \CM|dcif.imemload[8]~29_combout ;
wire \CM|dcif.imemload[7]~30_combout ;
wire \CM|dcif.imemload[6]~31_combout ;
wire \DP|ALU|Selector31~10_combout ;
wire \DP|ALU|ShiftRight0~50_combout ;
wire \DP|ALU|Selector24~0_combout ;
wire \DP|ALU|Selector8~0_combout ;
wire \DP|ALU|Selector0~33_combout ;
wire \DP|ALU|Selector3~10_combout ;
wire \DP|ALU|Selector4~1_combout ;
wire \DP|ALU|Selector7~17_combout ;
wire \DP|ALU|Selector11~8_combout ;
wire \DP|ALU|ShiftRight0~54_combout ;
wire \DP|ALU|Selector15~8_combout ;
wire \DP|ALU|Selector22~0_combout ;
wire \DP|ALU|Selector28~9_combout ;
wire \DP|ALU|Selector29~7_combout ;
wire \DP|ALU|ShiftRight0~85_combout ;
wire \DP|ALU|ShiftRight0~90_combout ;
wire \DP|ALU|ShiftLeft0~57_combout ;
wire \DP|ALU|Selector10~1_combout ;
wire \DP|ALU|Selector10~6_combout ;
wire \DP|ALU|Selector10~7_combout ;
wire \DP|ALU|Selector2~9_combout ;
wire \DP|ALU|Selector1~24_combout ;
wire \DP|ALU|Selector4~10_combout ;
wire \DP|ALU|Selector5~7_combout ;
wire \DP|ALU|Selector12~8_combout ;
wire \DP|ALU|Selector24~9_combout ;
wire \DP|ALU|Selector24~10_combout ;
wire \DP|ALU|Selector13~8_combout ;
wire \DP|ALU|Selector25~8_combout ;
wire \DP|ALU|Selector14~1_combout ;
wire \DP|ALU|Selector14~6_combout ;
wire \DP|ALU|Selector14~7_combout ;
wire \DP|ALU|Selector27~8_combout ;
wire \DP|ALU|Selector16~11_combout ;
wire \DP|ALU|Selector18~8_combout ;
wire \DP|ALU|Selector17~8_combout ;
wire \DP|ALU|Selector6~7_combout ;
wire \DP|ALU|Selector26~7_combout ;
wire \DP|ALU|Selector19~8_combout ;
wire \DP|ALU|Selector20~2_combout ;
wire \DP|ALU|Selector20~7_combout ;
wire \DP|ALU|Selector20~8_combout ;
wire \DP|ALU|Selector21~1_combout ;
wire \DP|ALU|Selector21~6_combout ;
wire \DP|ALU|Selector21~7_combout ;
wire \DP|ALU|Selector8~3_combout ;
wire \DP|ALU|Selector8~8_combout ;
wire \DP|ALU|Selector8~9_combout ;
wire \DP|ALU|Selector9~1_combout ;
wire \DP|ALU|Selector9~6_combout ;
wire \DP|ALU|Selector9~7_combout ;
wire \DP|ALU|Selector22~9_combout ;
wire \DP|ALU|Selector30~14_combout ;
wire \DP|ALU|Selector23~3_combout ;
wire \DP|ALU|Selector23~4_combout ;
wire \DP|ALU|Selector23~10_combout ;
wire \CM|dcif.dhit~0_combout ;
wire [31:0] \CM|instr ;


memory_control CC(
	.reg_WEN(reg_WEN),
	.reg_REN(reg_REN),
	.always1(always1),
	.ccifiwait_0(\CC|ccif.iwait[0]~0_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

caches CM(
	.daddr_1(daddr_1),
	.reg_WEN(reg_WEN),
	.reg_REN(reg_REN),
	.daddr_0(daddr_0),
	.daddr_3(daddr_3),
	.daddr_2(daddr_2),
	.daddr_5(daddr_5),
	.daddr_4(daddr_4),
	.daddr_7(daddr_7),
	.daddr_6(daddr_6),
	.daddr_9(daddr_9),
	.daddr_8(daddr_8),
	.daddr_11(daddr_11),
	.daddr_10(daddr_10),
	.daddr_13(daddr_13),
	.daddr_12(daddr_12),
	.daddr_15(daddr_15),
	.daddr_14(daddr_14),
	.daddr_17(daddr_17),
	.daddr_16(daddr_16),
	.daddr_19(daddr_19),
	.daddr_18(daddr_18),
	.daddr_21(daddr_21),
	.daddr_20(daddr_20),
	.daddr_23(daddr_23),
	.daddr_22(daddr_22),
	.daddr_25(daddr_25),
	.daddr_24(daddr_24),
	.daddr_27(daddr_27),
	.daddr_26(daddr_26),
	.daddr_29(daddr_29),
	.daddr_28(daddr_28),
	.daddr_31(daddr_31),
	.daddr_30(daddr_30),
	.always1(always1),
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.instr_30(\CM|instr [30]),
	.ccifiwait_0(\CC|ccif.iwait[0]~0_combout ),
	.dcifimemload_30(\CM|dcif.imemload[30]~0_combout ),
	.instr_31(\CM|instr [31]),
	.dcifimemload_31(\CM|dcif.imemload[31]~1_combout ),
	.instr_27(\CM|instr [27]),
	.dcifimemload_27(\CM|dcif.imemload[27]~2_combout ),
	.instr_26(\CM|instr [26]),
	.dcifimemload_26(\CM|dcif.imemload[26]~3_combout ),
	.instr_29(\CM|instr [29]),
	.dcifimemload_29(\CM|dcif.imemload[29]~4_combout ),
	.instr_28(\CM|instr [28]),
	.dcifimemload_28(\CM|dcif.imemload[28]~5_combout ),
	.dcifimemload_19(\CM|dcif.imemload[19]~6_combout ),
	.dcifimemload_18(\CM|dcif.imemload[18]~7_combout ),
	.instr_16(\CM|instr [16]),
	.dcifimemload_16(\CM|dcif.imemload[16]~8_combout ),
	.instr_17(\CM|instr [17]),
	.dcifimemload_17(\CM|dcif.imemload[17]~9_combout ),
	.dcifimemload_20(dcifimemload_20),
	.dcifimemload_24(\CM|dcif.imemload[24]~11_combout ),
	.dcifimemload_23(\CM|dcif.imemload[23]~12_combout ),
	.dcifimemload_21(\CM|dcif.imemload[21]~13_combout ),
	.dcifimemload_22(\CM|dcif.imemload[22]~14_combout ),
	.dcifimemload_25(\CM|dcif.imemload[25]~15_combout ),
	.dcifimemload_3(\CM|dcif.imemload[3]~16_combout ),
	.dcifimemload_4(\CM|dcif.imemload[4]~17_combout ),
	.dcifimemload_2(\CM|dcif.imemload[2]~18_combout ),
	.dcifimemload_5(\CM|dcif.imemload[5]~19_combout ),
	.dcifimemload_0(\CM|dcif.imemload[0]~20_combout ),
	.dcifimemload_1(\CM|dcif.imemload[1]~21_combout ),
	.dcifimemload_15(\CM|dcif.imemload[15]~22_combout ),
	.dcifimemload_14(\CM|dcif.imemload[14]~23_combout ),
	.dcifimemload_13(\CM|dcif.imemload[13]~24_combout ),
	.dcifimemload_12(\CM|dcif.imemload[12]~25_combout ),
	.dcifimemload_11(\CM|dcif.imemload[11]~26_combout ),
	.dcifimemload_10(\CM|dcif.imemload[10]~27_combout ),
	.dcifimemload_9(\CM|dcif.imemload[9]~28_combout ),
	.dcifimemload_8(\CM|dcif.imemload[8]~29_combout ),
	.dcifimemload_7(\CM|dcif.imemload[7]~30_combout ),
	.dcifimemload_6(\CM|dcif.imemload[6]~31_combout ),
	.Selector31(\DP|ALU|Selector31~10_combout ),
	.ShiftRight0(\DP|ALU|ShiftRight0~50_combout ),
	.Selector24(\DP|ALU|Selector24~0_combout ),
	.Selector8(\DP|ALU|Selector8~0_combout ),
	.Selector0(\DP|ALU|Selector0~33_combout ),
	.Selector3(\DP|ALU|Selector3~10_combout ),
	.Selector4(\DP|ALU|Selector4~1_combout ),
	.Selector7(\DP|ALU|Selector7~17_combout ),
	.Selector11(\DP|ALU|Selector11~8_combout ),
	.ShiftRight01(\DP|ALU|ShiftRight0~54_combout ),
	.Selector15(\DP|ALU|Selector15~8_combout ),
	.Selector22(\DP|ALU|Selector22~0_combout ),
	.Selector28(\DP|ALU|Selector28~9_combout ),
	.Selector29(\DP|ALU|Selector29~7_combout ),
	.ShiftRight02(\DP|ALU|ShiftRight0~85_combout ),
	.ShiftRight03(\DP|ALU|ShiftRight0~90_combout ),
	.ShiftLeft0(\DP|ALU|ShiftLeft0~57_combout ),
	.Selector10(\DP|ALU|Selector10~1_combout ),
	.Selector101(\DP|ALU|Selector10~6_combout ),
	.Selector102(\DP|ALU|Selector10~7_combout ),
	.Selector2(\DP|ALU|Selector2~9_combout ),
	.Selector1(\DP|ALU|Selector1~24_combout ),
	.Selector41(\DP|ALU|Selector4~10_combout ),
	.Selector5(\DP|ALU|Selector5~7_combout ),
	.Selector12(\DP|ALU|Selector12~8_combout ),
	.Selector241(\DP|ALU|Selector24~9_combout ),
	.Selector242(\DP|ALU|Selector24~10_combout ),
	.Selector13(\DP|ALU|Selector13~8_combout ),
	.Selector25(\DP|ALU|Selector25~8_combout ),
	.Selector14(\DP|ALU|Selector14~1_combout ),
	.Selector141(\DP|ALU|Selector14~6_combout ),
	.Selector142(\DP|ALU|Selector14~7_combout ),
	.Selector27(\DP|ALU|Selector27~8_combout ),
	.Selector16(\DP|ALU|Selector16~11_combout ),
	.Selector18(\DP|ALU|Selector18~8_combout ),
	.Selector17(\DP|ALU|Selector17~8_combout ),
	.Selector6(\DP|ALU|Selector6~7_combout ),
	.Selector26(\DP|ALU|Selector26~7_combout ),
	.Selector19(\DP|ALU|Selector19~8_combout ),
	.Selector20(\DP|ALU|Selector20~2_combout ),
	.Selector201(\DP|ALU|Selector20~7_combout ),
	.Selector202(\DP|ALU|Selector20~8_combout ),
	.Selector21(\DP|ALU|Selector21~1_combout ),
	.Selector211(\DP|ALU|Selector21~6_combout ),
	.Selector212(\DP|ALU|Selector21~7_combout ),
	.Selector81(\DP|ALU|Selector8~3_combout ),
	.Selector82(\DP|ALU|Selector8~8_combout ),
	.Selector83(\DP|ALU|Selector8~9_combout ),
	.Selector9(\DP|ALU|Selector9~1_combout ),
	.Selector91(\DP|ALU|Selector9~6_combout ),
	.Selector92(\DP|ALU|Selector9~7_combout ),
	.Selector221(\DP|ALU|Selector22~9_combout ),
	.Selector30(\DP|ALU|Selector30~14_combout ),
	.Selector23(\DP|ALU|Selector23~3_combout ),
	.Selector231(\DP|ALU|Selector23~4_combout ),
	.Selector232(\DP|ALU|Selector23~10_combout ),
	.dcifdhit(\CM|dcif.dhit~0_combout ),
	.nRST(nRST),
	.CLK(CLK),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

datapath DP(
	.PC_29(PC_29),
	.PC_28(PC_28),
	.PC_31(PC_31),
	.PC_30(PC_30),
	.dpifhalt(dpifhalt),
	.PC_1(PC_1),
	.reg_WEN(reg_WEN),
	.reg_REN(reg_REN),
	.PC_0(PC_0),
	.PC_3(PC_3),
	.PC_2(PC_2),
	.PC_5(PC_5),
	.PC_4(PC_4),
	.PC_7(PC_7),
	.PC_6(PC_6),
	.PC_9(PC_9),
	.PC_8(PC_8),
	.PC_11(PC_11),
	.PC_10(PC_10),
	.PC_13(PC_13),
	.PC_12(PC_12),
	.PC_15(PC_15),
	.PC_14(PC_14),
	.PC_17(PC_17),
	.PC_16(PC_16),
	.PC_19(PC_19),
	.PC_18(PC_18),
	.PC_21(PC_21),
	.PC_20(PC_20),
	.PC_23(PC_23),
	.PC_22(PC_22),
	.PC_25(PC_25),
	.PC_24(PC_24),
	.PC_27(PC_27),
	.PC_26(PC_26),
	.always1(always1),
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.instr_30(\CM|instr [30]),
	.ccifiwait_0(\CC|ccif.iwait[0]~0_combout ),
	.dcifimemload_30(\CM|dcif.imemload[30]~0_combout ),
	.instr_31(\CM|instr [31]),
	.dcifimemload_31(\CM|dcif.imemload[31]~1_combout ),
	.instr_27(\CM|instr [27]),
	.dcifimemload_27(\CM|dcif.imemload[27]~2_combout ),
	.instr_26(\CM|instr [26]),
	.dcifimemload_26(\CM|dcif.imemload[26]~3_combout ),
	.instr_29(\CM|instr [29]),
	.dcifimemload_29(\CM|dcif.imemload[29]~4_combout ),
	.instr_28(\CM|instr [28]),
	.dcifimemload_28(\CM|dcif.imemload[28]~5_combout ),
	.dcifimemload_19(\CM|dcif.imemload[19]~6_combout ),
	.dcifimemload_18(\CM|dcif.imemload[18]~7_combout ),
	.instr_16(\CM|instr [16]),
	.dcifimemload_16(\CM|dcif.imemload[16]~8_combout ),
	.instr_17(\CM|instr [17]),
	.dcifimemload_17(\CM|dcif.imemload[17]~9_combout ),
	.Mux63(Mux63),
	.Mux631(Mux631),
	.dcifimemload_20(dcifimemload_20),
	.dcifimemload_24(\CM|dcif.imemload[24]~11_combout ),
	.dcifimemload_23(\CM|dcif.imemload[23]~12_combout ),
	.dcifimemload_21(\CM|dcif.imemload[21]~13_combout ),
	.dcifimemload_22(\CM|dcif.imemload[22]~14_combout ),
	.dcifimemload_25(\CM|dcif.imemload[25]~15_combout ),
	.dcifimemload_3(\CM|dcif.imemload[3]~16_combout ),
	.dcifimemload_4(\CM|dcif.imemload[4]~17_combout ),
	.dcifimemload_2(\CM|dcif.imemload[2]~18_combout ),
	.dcifimemload_5(\CM|dcif.imemload[5]~19_combout ),
	.dcifimemload_0(\CM|dcif.imemload[0]~20_combout ),
	.dcifimemload_1(\CM|dcif.imemload[1]~21_combout ),
	.dcifimemload_15(\CM|dcif.imemload[15]~22_combout ),
	.Mux32(Mux32),
	.Mux321(Mux321),
	.Mux33(Mux33),
	.Mux331(Mux331),
	.Mux34(Mux34),
	.Mux341(Mux341),
	.Mux35(Mux35),
	.Mux351(Mux351),
	.Mux36(Mux36),
	.Mux361(Mux361),
	.Mux37(Mux37),
	.Mux371(Mux371),
	.Mux38(Mux38),
	.Mux381(Mux381),
	.Mux39(Mux39),
	.Mux391(Mux391),
	.Mux40(Mux40),
	.Mux401(Mux401),
	.Mux41(Mux41),
	.Mux411(Mux411),
	.Mux42(Mux42),
	.Mux421(Mux421),
	.Mux43(Mux43),
	.Mux431(Mux431),
	.Mux44(Mux44),
	.Mux441(Mux441),
	.Mux45(Mux45),
	.Mux451(Mux451),
	.Mux46(Mux46),
	.Mux461(Mux461),
	.Mux47(Mux47),
	.Mux471(Mux471),
	.Mux48(Mux48),
	.Mux481(Mux481),
	.dcifimemload_14(\CM|dcif.imemload[14]~23_combout ),
	.Mux49(Mux49),
	.Mux491(Mux491),
	.dcifimemload_13(\CM|dcif.imemload[13]~24_combout ),
	.Mux50(Mux50),
	.Mux501(Mux501),
	.dcifimemload_12(\CM|dcif.imemload[12]~25_combout ),
	.Mux51(Mux51),
	.Mux511(Mux511),
	.dcifimemload_11(\CM|dcif.imemload[11]~26_combout ),
	.Mux52(Mux52),
	.Mux521(Mux521),
	.dcifimemload_10(\CM|dcif.imemload[10]~27_combout ),
	.Mux53(Mux53),
	.Mux531(Mux531),
	.dcifimemload_9(\CM|dcif.imemload[9]~28_combout ),
	.Mux54(Mux54),
	.Mux541(Mux541),
	.dcifimemload_8(\CM|dcif.imemload[8]~29_combout ),
	.Mux55(Mux55),
	.Mux551(Mux551),
	.dcifimemload_7(\CM|dcif.imemload[7]~30_combout ),
	.Mux56(Mux56),
	.Mux561(Mux561),
	.dcifimemload_6(\CM|dcif.imemload[6]~31_combout ),
	.Mux57(Mux57),
	.Mux571(Mux571),
	.Mux58(Mux58),
	.Mux581(Mux581),
	.Mux59(Mux59),
	.Mux591(Mux591),
	.Mux60(Mux60),
	.Mux601(Mux601),
	.Mux61(Mux61),
	.Mux611(Mux611),
	.Mux62(Mux62),
	.Mux621(Mux621),
	.Selector31(\DP|ALU|Selector31~10_combout ),
	.ShiftRight0(\DP|ALU|ShiftRight0~50_combout ),
	.Selector24(\DP|ALU|Selector24~0_combout ),
	.Selector8(\DP|ALU|Selector8~0_combout ),
	.Selector0(\DP|ALU|Selector0~33_combout ),
	.Selector3(\DP|ALU|Selector3~10_combout ),
	.Selector4(\DP|ALU|Selector4~1_combout ),
	.Selector7(\DP|ALU|Selector7~17_combout ),
	.Selector11(\DP|ALU|Selector11~8_combout ),
	.ShiftRight01(\DP|ALU|ShiftRight0~54_combout ),
	.Selector15(\DP|ALU|Selector15~8_combout ),
	.Selector22(\DP|ALU|Selector22~0_combout ),
	.Selector28(\DP|ALU|Selector28~9_combout ),
	.Selector29(\DP|ALU|Selector29~7_combout ),
	.ShiftRight02(\DP|ALU|ShiftRight0~85_combout ),
	.ShiftRight03(\DP|ALU|ShiftRight0~90_combout ),
	.ShiftLeft0(\DP|ALU|ShiftLeft0~57_combout ),
	.Selector10(\DP|ALU|Selector10~1_combout ),
	.Selector101(\DP|ALU|Selector10~6_combout ),
	.Selector102(\DP|ALU|Selector10~7_combout ),
	.Selector2(\DP|ALU|Selector2~9_combout ),
	.Selector1(\DP|ALU|Selector1~24_combout ),
	.Selector41(\DP|ALU|Selector4~10_combout ),
	.Selector5(\DP|ALU|Selector5~7_combout ),
	.Selector12(\DP|ALU|Selector12~8_combout ),
	.Selector241(\DP|ALU|Selector24~9_combout ),
	.Selector242(\DP|ALU|Selector24~10_combout ),
	.Selector13(\DP|ALU|Selector13~8_combout ),
	.Selector25(\DP|ALU|Selector25~8_combout ),
	.Selector14(\DP|ALU|Selector14~1_combout ),
	.Selector141(\DP|ALU|Selector14~6_combout ),
	.Selector142(\DP|ALU|Selector14~7_combout ),
	.Selector27(\DP|ALU|Selector27~8_combout ),
	.Selector16(\DP|ALU|Selector16~11_combout ),
	.Selector18(\DP|ALU|Selector18~8_combout ),
	.Selector17(\DP|ALU|Selector17~8_combout ),
	.Selector6(\DP|ALU|Selector6~7_combout ),
	.Selector26(\DP|ALU|Selector26~7_combout ),
	.Selector19(\DP|ALU|Selector19~8_combout ),
	.Selector20(\DP|ALU|Selector20~2_combout ),
	.Selector201(\DP|ALU|Selector20~7_combout ),
	.Selector202(\DP|ALU|Selector20~8_combout ),
	.Selector21(\DP|ALU|Selector21~1_combout ),
	.Selector211(\DP|ALU|Selector21~6_combout ),
	.Selector212(\DP|ALU|Selector21~7_combout ),
	.Selector81(\DP|ALU|Selector8~3_combout ),
	.Selector82(\DP|ALU|Selector8~8_combout ),
	.Selector83(\DP|ALU|Selector8~9_combout ),
	.Selector9(\DP|ALU|Selector9~1_combout ),
	.Selector91(\DP|ALU|Selector9~6_combout ),
	.Selector92(\DP|ALU|Selector9~7_combout ),
	.Selector221(\DP|ALU|Selector22~9_combout ),
	.Selector30(\DP|ALU|Selector30~14_combout ),
	.Selector23(\DP|ALU|Selector23~3_combout ),
	.Selector231(\DP|ALU|Selector23~4_combout ),
	.Selector232(\DP|ALU|Selector23~10_combout ),
	.dcifdhit(\CM|dcif.dhit~0_combout ),
	.CLK(CLK),
	.nRST(nRST1),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module caches (
	daddr_1,
	reg_WEN,
	reg_REN,
	daddr_0,
	daddr_3,
	daddr_2,
	daddr_5,
	daddr_4,
	daddr_7,
	daddr_6,
	daddr_9,
	daddr_8,
	daddr_11,
	daddr_10,
	daddr_13,
	daddr_12,
	daddr_15,
	daddr_14,
	daddr_17,
	daddr_16,
	daddr_19,
	daddr_18,
	daddr_21,
	daddr_20,
	daddr_23,
	daddr_22,
	daddr_25,
	daddr_24,
	daddr_27,
	daddr_26,
	daddr_29,
	daddr_28,
	daddr_31,
	daddr_30,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	instr_30,
	ccifiwait_0,
	dcifimemload_30,
	instr_31,
	dcifimemload_31,
	instr_27,
	dcifimemload_27,
	instr_26,
	dcifimemload_26,
	instr_29,
	dcifimemload_29,
	instr_28,
	dcifimemload_28,
	dcifimemload_19,
	dcifimemload_18,
	instr_16,
	dcifimemload_16,
	instr_17,
	dcifimemload_17,
	dcifimemload_20,
	dcifimemload_24,
	dcifimemload_23,
	dcifimemload_21,
	dcifimemload_22,
	dcifimemload_25,
	dcifimemload_3,
	dcifimemload_4,
	dcifimemload_2,
	dcifimemload_5,
	dcifimemload_0,
	dcifimemload_1,
	dcifimemload_15,
	dcifimemload_14,
	dcifimemload_13,
	dcifimemload_12,
	dcifimemload_11,
	dcifimemload_10,
	dcifimemload_9,
	dcifimemload_8,
	dcifimemload_7,
	dcifimemload_6,
	Selector31,
	ShiftRight0,
	Selector24,
	Selector8,
	Selector0,
	Selector3,
	Selector4,
	Selector7,
	Selector11,
	ShiftRight01,
	Selector15,
	Selector22,
	Selector28,
	Selector29,
	ShiftRight02,
	ShiftRight03,
	ShiftLeft0,
	Selector10,
	Selector101,
	Selector102,
	Selector2,
	Selector1,
	Selector41,
	Selector5,
	Selector12,
	Selector241,
	Selector242,
	Selector13,
	Selector25,
	Selector14,
	Selector141,
	Selector142,
	Selector27,
	Selector16,
	Selector18,
	Selector17,
	Selector6,
	Selector26,
	Selector19,
	Selector20,
	Selector201,
	Selector202,
	Selector21,
	Selector211,
	Selector212,
	Selector81,
	Selector82,
	Selector83,
	Selector9,
	Selector91,
	Selector92,
	Selector221,
	Selector30,
	Selector23,
	Selector231,
	Selector232,
	dcifdhit,
	nRST,
	CLK,
	devpor,
	devclrn,
	devoe);
output 	daddr_1;
input 	reg_WEN;
input 	reg_REN;
output 	daddr_0;
output 	daddr_3;
output 	daddr_2;
output 	daddr_5;
output 	daddr_4;
output 	daddr_7;
output 	daddr_6;
output 	daddr_9;
output 	daddr_8;
output 	daddr_11;
output 	daddr_10;
output 	daddr_13;
output 	daddr_12;
output 	daddr_15;
output 	daddr_14;
output 	daddr_17;
output 	daddr_16;
output 	daddr_19;
output 	daddr_18;
output 	daddr_21;
output 	daddr_20;
output 	daddr_23;
output 	daddr_22;
output 	daddr_25;
output 	daddr_24;
output 	daddr_27;
output 	daddr_26;
output 	daddr_29;
output 	daddr_28;
output 	daddr_31;
output 	daddr_30;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
output 	instr_30;
input 	ccifiwait_0;
output 	dcifimemload_30;
output 	instr_31;
output 	dcifimemload_31;
output 	instr_27;
output 	dcifimemload_27;
output 	instr_26;
output 	dcifimemload_26;
output 	instr_29;
output 	dcifimemload_29;
output 	instr_28;
output 	dcifimemload_28;
output 	dcifimemload_19;
output 	dcifimemload_18;
output 	instr_16;
output 	dcifimemload_16;
output 	instr_17;
output 	dcifimemload_17;
output 	dcifimemload_20;
output 	dcifimemload_24;
output 	dcifimemload_23;
output 	dcifimemload_21;
output 	dcifimemload_22;
output 	dcifimemload_25;
output 	dcifimemload_3;
output 	dcifimemload_4;
output 	dcifimemload_2;
output 	dcifimemload_5;
output 	dcifimemload_0;
output 	dcifimemload_1;
output 	dcifimemload_15;
output 	dcifimemload_14;
output 	dcifimemload_13;
output 	dcifimemload_12;
output 	dcifimemload_11;
output 	dcifimemload_10;
output 	dcifimemload_9;
output 	dcifimemload_8;
output 	dcifimemload_7;
output 	dcifimemload_6;
input 	Selector31;
input 	ShiftRight0;
input 	Selector24;
input 	Selector8;
input 	Selector0;
input 	Selector3;
input 	Selector4;
input 	Selector7;
input 	Selector11;
input 	ShiftRight01;
input 	Selector15;
input 	Selector22;
input 	Selector28;
input 	Selector29;
input 	ShiftRight02;
input 	ShiftRight03;
input 	ShiftLeft0;
input 	Selector10;
input 	Selector101;
input 	Selector102;
input 	Selector2;
input 	Selector1;
input 	Selector41;
input 	Selector5;
input 	Selector12;
input 	Selector241;
input 	Selector242;
input 	Selector13;
input 	Selector25;
input 	Selector14;
input 	Selector141;
input 	Selector142;
input 	Selector27;
input 	Selector16;
input 	Selector18;
input 	Selector17;
input 	Selector6;
input 	Selector26;
input 	Selector19;
input 	Selector20;
input 	Selector201;
input 	Selector202;
input 	Selector21;
input 	Selector211;
input 	Selector212;
input 	Selector81;
input 	Selector82;
input 	Selector83;
input 	Selector9;
input 	Selector91;
input 	Selector92;
input 	Selector221;
input 	Selector30;
input 	Selector23;
input 	Selector231;
input 	Selector232;
output 	dcifdhit;
input 	nRST;
input 	CLK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \daddr~0_combout ;
wire \daddr[1]~1_combout ;
wire \daddr~2_combout ;
wire \daddr~3_combout ;
wire \daddr~4_combout ;
wire \daddr~5_combout ;
wire \daddr~6_combout ;
wire \daddr~7_combout ;
wire \daddr~8_combout ;
wire \daddr~9_combout ;
wire \daddr~10_combout ;
wire \daddr~11_combout ;
wire \daddr~12_combout ;
wire \daddr~13_combout ;
wire \daddr~14_combout ;
wire \daddr~15_combout ;
wire \daddr~16_combout ;
wire \daddr~17_combout ;
wire \daddr~18_combout ;
wire \daddr~19_combout ;
wire \daddr~20_combout ;
wire \daddr~21_combout ;
wire \daddr~22_combout ;
wire \daddr~23_combout ;
wire \daddr~24_combout ;
wire \daddr~25_combout ;
wire \daddr~26_combout ;
wire \daddr~27_combout ;
wire \daddr~28_combout ;
wire \daddr~29_combout ;
wire \daddr~30_combout ;
wire \daddr~31_combout ;
wire \daddr~32_combout ;
wire \instr~0_combout ;
wire \instr~1_combout ;
wire \instr~2_combout ;
wire \instr~3_combout ;
wire \instr~4_combout ;
wire \instr~5_combout ;
wire \instr~6_combout ;
wire \instr~7_combout ;
wire \instr~8_combout ;
wire \instr[16]~feeder_combout ;
wire \instr~9_combout ;
wire \instr~10_combout ;
wire \instr~11_combout ;
wire \instr~12_combout ;
wire \instr~13_combout ;
wire \instr~14_combout ;
wire \instr~15_combout ;
wire \instr~16_combout ;
wire \instr~17_combout ;
wire \instr~18_combout ;
wire \instr~19_combout ;
wire \instr~20_combout ;
wire \instr~21_combout ;
wire \instr~22_combout ;
wire \instr~23_combout ;
wire \instr~24_combout ;
wire \instr~25_combout ;
wire \instr~26_combout ;
wire \instr~27_combout ;
wire \instr~28_combout ;
wire \instr~29_combout ;
wire \instr~30_combout ;
wire \instr~31_combout ;
wire [31:0] instr;


// Location: FF_X60_Y33_N25
dffeas \daddr[1] (
	.clk(CLK),
	.d(\daddr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_1),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[1] .is_wysiwyg = "true";
defparam \daddr[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N27
dffeas \daddr[0] (
	.clk(CLK),
	.d(\daddr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_0),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[0] .is_wysiwyg = "true";
defparam \daddr[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N13
dffeas \daddr[3] (
	.clk(CLK),
	.d(\daddr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_3),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[3] .is_wysiwyg = "true";
defparam \daddr[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N31
dffeas \daddr[2] (
	.clk(CLK),
	.d(\daddr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_2),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[2] .is_wysiwyg = "true";
defparam \daddr[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N23
dffeas \daddr[5] (
	.clk(CLK),
	.d(\daddr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_5),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[5] .is_wysiwyg = "true";
defparam \daddr[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N1
dffeas \daddr[4] (
	.clk(CLK),
	.d(\daddr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_4),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[4] .is_wysiwyg = "true";
defparam \daddr[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N5
dffeas \daddr[7] (
	.clk(CLK),
	.d(\daddr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_7),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[7] .is_wysiwyg = "true";
defparam \daddr[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N27
dffeas \daddr[6] (
	.clk(CLK),
	.d(\daddr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_6),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[6] .is_wysiwyg = "true";
defparam \daddr[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N29
dffeas \daddr[9] (
	.clk(CLK),
	.d(\daddr~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_9),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[9] .is_wysiwyg = "true";
defparam \daddr[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N15
dffeas \daddr[8] (
	.clk(CLK),
	.d(\daddr~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_8),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[8] .is_wysiwyg = "true";
defparam \daddr[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N13
dffeas \daddr[11] (
	.clk(CLK),
	.d(\daddr~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_11),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[11] .is_wysiwyg = "true";
defparam \daddr[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N25
dffeas \daddr[10] (
	.clk(CLK),
	.d(\daddr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_10),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[10] .is_wysiwyg = "true";
defparam \daddr[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y35_N21
dffeas \daddr[13] (
	.clk(CLK),
	.d(\daddr~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_13),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[13] .is_wysiwyg = "true";
defparam \daddr[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y35_N15
dffeas \daddr[12] (
	.clk(CLK),
	.d(\daddr~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_12),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[12] .is_wysiwyg = "true";
defparam \daddr[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N29
dffeas \daddr[15] (
	.clk(CLK),
	.d(\daddr~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_15),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[15] .is_wysiwyg = "true";
defparam \daddr[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N31
dffeas \daddr[14] (
	.clk(CLK),
	.d(\daddr~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_14),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[14] .is_wysiwyg = "true";
defparam \daddr[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N3
dffeas \daddr[17] (
	.clk(CLK),
	.d(\daddr~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_17),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[17] .is_wysiwyg = "true";
defparam \daddr[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y34_N5
dffeas \daddr[16] (
	.clk(CLK),
	.d(\daddr~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_16),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[16] .is_wysiwyg = "true";
defparam \daddr[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N17
dffeas \daddr[19] (
	.clk(CLK),
	.d(\daddr~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_19),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[19] .is_wysiwyg = "true";
defparam \daddr[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N25
dffeas \daddr[18] (
	.clk(CLK),
	.d(\daddr~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_18),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[18] .is_wysiwyg = "true";
defparam \daddr[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N5
dffeas \daddr[21] (
	.clk(CLK),
	.d(\daddr~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_21),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[21] .is_wysiwyg = "true";
defparam \daddr[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N31
dffeas \daddr[20] (
	.clk(CLK),
	.d(\daddr~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_20),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[20] .is_wysiwyg = "true";
defparam \daddr[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N15
dffeas \daddr[23] (
	.clk(CLK),
	.d(\daddr~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_23),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[23] .is_wysiwyg = "true";
defparam \daddr[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N5
dffeas \daddr[22] (
	.clk(CLK),
	.d(\daddr~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_22),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[22] .is_wysiwyg = "true";
defparam \daddr[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N5
dffeas \daddr[25] (
	.clk(CLK),
	.d(\daddr~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_25),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[25] .is_wysiwyg = "true";
defparam \daddr[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N27
dffeas \daddr[24] (
	.clk(CLK),
	.d(\daddr~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_24),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[24] .is_wysiwyg = "true";
defparam \daddr[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N29
dffeas \daddr[27] (
	.clk(CLK),
	.d(\daddr~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_27),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[27] .is_wysiwyg = "true";
defparam \daddr[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N5
dffeas \daddr[26] (
	.clk(CLK),
	.d(\daddr~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_26),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[26] .is_wysiwyg = "true";
defparam \daddr[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N25
dffeas \daddr[29] (
	.clk(CLK),
	.d(\daddr~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_29),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[29] .is_wysiwyg = "true";
defparam \daddr[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N13
dffeas \daddr[28] (
	.clk(CLK),
	.d(\daddr~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_28),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[28] .is_wysiwyg = "true";
defparam \daddr[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N17
dffeas \daddr[31] (
	.clk(CLK),
	.d(\daddr~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_31),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[31] .is_wysiwyg = "true";
defparam \daddr[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N9
dffeas \daddr[30] (
	.clk(CLK),
	.d(\daddr~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_30),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[30] .is_wysiwyg = "true";
defparam \daddr[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y30_N5
dffeas \instr[30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~0_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_30),
	.prn(vcc));
// synopsys translate_off
defparam \instr[30] .is_wysiwyg = "true";
defparam \instr[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N10
cycloneive_lcell_comb \dcif.imemload[30]~0 (
// Equation(s):
// dcifimemload_30 = (ccifiwait_0 & ((ramiframload_30))) # (!ccifiwait_0 & (instr_30))

	.dataa(gnd),
	.datab(instr_30),
	.datac(ramiframload_30),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_30),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[30]~0 .lut_mask = 16'hF0CC;
defparam \dcif.imemload[30]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y30_N21
dffeas \instr[31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_31),
	.prn(vcc));
// synopsys translate_off
defparam \instr[31] .is_wysiwyg = "true";
defparam \instr[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N20
cycloneive_lcell_comb \dcif.imemload[31]~1 (
// Equation(s):
// dcifimemload_31 = (ccifiwait_0 & (ramiframload_31)) # (!ccifiwait_0 & ((instr_31)))

	.dataa(gnd),
	.datab(ramiframload_31),
	.datac(instr_31),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_31),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[31]~1 .lut_mask = 16'hCCF0;
defparam \dcif.imemload[31]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y30_N19
dffeas \instr[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_27),
	.prn(vcc));
// synopsys translate_off
defparam \instr[27] .is_wysiwyg = "true";
defparam \instr[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N20
cycloneive_lcell_comb \dcif.imemload[27]~2 (
// Equation(s):
// dcifimemload_27 = (ccifiwait_0 & ((ramiframload_27))) # (!ccifiwait_0 & (instr_27))

	.dataa(gnd),
	.datab(instr_27),
	.datac(ccifiwait_0),
	.datad(ramiframload_27),
	.cin(gnd),
	.combout(dcifimemload_27),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[27]~2 .lut_mask = 16'hFC0C;
defparam \dcif.imemload[27]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y30_N23
dffeas \instr[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_26),
	.prn(vcc));
// synopsys translate_off
defparam \instr[26] .is_wysiwyg = "true";
defparam \instr[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N12
cycloneive_lcell_comb \dcif.imemload[26]~3 (
// Equation(s):
// dcifimemload_26 = (ccifiwait_0 & ((ramiframload_26))) # (!ccifiwait_0 & (instr_26))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr_26),
	.datad(ramiframload_26),
	.cin(gnd),
	.combout(dcifimemload_26),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[26]~3 .lut_mask = 16'hFC30;
defparam \dcif.imemload[26]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y30_N21
dffeas \instr[29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_29),
	.prn(vcc));
// synopsys translate_off
defparam \instr[29] .is_wysiwyg = "true";
defparam \instr[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N20
cycloneive_lcell_comb \dcif.imemload[29]~4 (
// Equation(s):
// dcifimemload_29 = (ccifiwait_0 & ((ramiframload_29))) # (!ccifiwait_0 & (instr_29))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(instr_29),
	.datad(ramiframload_29),
	.cin(gnd),
	.combout(dcifimemload_29),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[29]~4 .lut_mask = 16'hFA50;
defparam \dcif.imemload[29]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N25
dffeas \instr[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_28),
	.prn(vcc));
// synopsys translate_off
defparam \instr[28] .is_wysiwyg = "true";
defparam \instr[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N22
cycloneive_lcell_comb \dcif.imemload[28]~5 (
// Equation(s):
// dcifimemload_28 = (ccifiwait_0 & ((ramiframload_28))) # (!ccifiwait_0 & (instr_28))

	.dataa(gnd),
	.datab(instr_28),
	.datac(ramiframload_28),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_28),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[28]~5 .lut_mask = 16'hF0CC;
defparam \dcif.imemload[28]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N20
cycloneive_lcell_comb \dcif.imemload[19]~6 (
// Equation(s):
// dcifimemload_19 = (ccifiwait_0 & (ramiframload_19)) # (!ccifiwait_0 & ((instr[19])))

	.dataa(ramiframload_19),
	.datab(gnd),
	.datac(instr[19]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_19),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[19]~6 .lut_mask = 16'hAAF0;
defparam \dcif.imemload[19]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N28
cycloneive_lcell_comb \dcif.imemload[18]~7 (
// Equation(s):
// dcifimemload_18 = (ccifiwait_0 & (ramiframload_18)) # (!ccifiwait_0 & ((instr[18])))

	.dataa(ramiframload_18),
	.datab(gnd),
	.datac(instr[18]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_18),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[18]~7 .lut_mask = 16'hAAF0;
defparam \dcif.imemload[18]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N25
dffeas \instr[16] (
	.clk(CLK),
	.d(\instr[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_16),
	.prn(vcc));
// synopsys translate_off
defparam \instr[16] .is_wysiwyg = "true";
defparam \instr[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N6
cycloneive_lcell_comb \dcif.imemload[16]~8 (
// Equation(s):
// dcifimemload_16 = (ccifiwait_0 & ((ramiframload_16))) # (!ccifiwait_0 & (instr_16))

	.dataa(gnd),
	.datab(instr_16),
	.datac(ccifiwait_0),
	.datad(ramiframload_16),
	.cin(gnd),
	.combout(dcifimemload_16),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[16]~8 .lut_mask = 16'hFC0C;
defparam \dcif.imemload[16]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N17
dffeas \instr[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~9_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_17),
	.prn(vcc));
// synopsys translate_off
defparam \instr[17] .is_wysiwyg = "true";
defparam \instr[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N2
cycloneive_lcell_comb \dcif.imemload[17]~9 (
// Equation(s):
// dcifimemload_17 = (ccifiwait_0 & ((ramiframload_17))) # (!ccifiwait_0 & (instr_17))

	.dataa(gnd),
	.datab(instr_17),
	.datac(ccifiwait_0),
	.datad(ramiframload_17),
	.cin(gnd),
	.combout(dcifimemload_17),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[17]~9 .lut_mask = 16'hFC0C;
defparam \dcif.imemload[17]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N18
cycloneive_lcell_comb \dcif.imemload[20]~10 (
// Equation(s):
// dcifimemload_20 = (ccifiwait_0 & (ramiframload_20)) # (!ccifiwait_0 & ((instr[20])))

	.dataa(gnd),
	.datab(ramiframload_20),
	.datac(instr[20]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_20),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[20]~10 .lut_mask = 16'hCCF0;
defparam \dcif.imemload[20]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N14
cycloneive_lcell_comb \dcif.imemload[24]~11 (
// Equation(s):
// dcifimemload_24 = (ccifiwait_0 & ((ramiframload_24))) # (!ccifiwait_0 & (instr[24]))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[24]),
	.datad(ramiframload_24),
	.cin(gnd),
	.combout(dcifimemload_24),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[24]~11 .lut_mask = 16'hFC30;
defparam \dcif.imemload[24]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N0
cycloneive_lcell_comb \dcif.imemload[23]~12 (
// Equation(s):
// dcifimemload_23 = (ccifiwait_0 & ((ramiframload_23))) # (!ccifiwait_0 & (instr[23]))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[23]),
	.datad(ramiframload_23),
	.cin(gnd),
	.combout(dcifimemload_23),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[23]~12 .lut_mask = 16'hFC30;
defparam \dcif.imemload[23]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N0
cycloneive_lcell_comb \dcif.imemload[21]~13 (
// Equation(s):
// dcifimemload_21 = (ccifiwait_0 & (ramiframload_21)) # (!ccifiwait_0 & ((instr[21])))

	.dataa(ramiframload_21),
	.datab(gnd),
	.datac(instr[21]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_21),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[21]~13 .lut_mask = 16'hAAF0;
defparam \dcif.imemload[21]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N16
cycloneive_lcell_comb \dcif.imemload[22]~14 (
// Equation(s):
// dcifimemload_22 = (ccifiwait_0 & (ramiframload_22)) # (!ccifiwait_0 & ((instr[22])))

	.dataa(gnd),
	.datab(ramiframload_22),
	.datac(instr[22]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_22),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[22]~14 .lut_mask = 16'hCCF0;
defparam \dcif.imemload[22]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N10
cycloneive_lcell_comb \dcif.imemload[25]~15 (
// Equation(s):
// dcifimemload_25 = (ccifiwait_0 & (ramiframload_25)) # (!ccifiwait_0 & ((instr[25])))

	.dataa(gnd),
	.datab(ramiframload_25),
	.datac(instr[25]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_25),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[25]~15 .lut_mask = 16'hCCF0;
defparam \dcif.imemload[25]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N0
cycloneive_lcell_comb \dcif.imemload[3]~16 (
// Equation(s):
// dcifimemload_3 = (ccifiwait_0 & (ramiframload_3)) # (!ccifiwait_0 & ((instr[3])))

	.dataa(gnd),
	.datab(ramiframload_3),
	.datac(instr[3]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_3),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[3]~16 .lut_mask = 16'hCCF0;
defparam \dcif.imemload[3]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N24
cycloneive_lcell_comb \dcif.imemload[4]~17 (
// Equation(s):
// dcifimemload_4 = (ccifiwait_0 & ((ramiframload_4))) # (!ccifiwait_0 & (instr[4]))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(instr[4]),
	.datad(ramiframload_4),
	.cin(gnd),
	.combout(dcifimemload_4),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[4]~17 .lut_mask = 16'hFA50;
defparam \dcif.imemload[4]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N30
cycloneive_lcell_comb \dcif.imemload[2]~18 (
// Equation(s):
// dcifimemload_2 = (ccifiwait_0 & (ramiframload_2)) # (!ccifiwait_0 & ((instr[2])))

	.dataa(ramiframload_2),
	.datab(gnd),
	.datac(instr[2]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_2),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[2]~18 .lut_mask = 16'hAAF0;
defparam \dcif.imemload[2]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N16
cycloneive_lcell_comb \dcif.imemload[5]~19 (
// Equation(s):
// dcifimemload_5 = (ccifiwait_0 & (ramiframload_5)) # (!ccifiwait_0 & ((instr[5])))

	.dataa(gnd),
	.datab(ramiframload_5),
	.datac(instr[5]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_5),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[5]~19 .lut_mask = 16'hCCF0;
defparam \dcif.imemload[5]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N30
cycloneive_lcell_comb \dcif.imemload[0]~20 (
// Equation(s):
// dcifimemload_0 = (ccifiwait_0 & ((ramiframload_0))) # (!ccifiwait_0 & (instr[0]))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(instr[0]),
	.datad(ramiframload_0),
	.cin(gnd),
	.combout(dcifimemload_0),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[0]~20 .lut_mask = 16'hFA50;
defparam \dcif.imemload[0]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N28
cycloneive_lcell_comb \dcif.imemload[1]~21 (
// Equation(s):
// dcifimemload_1 = (ccifiwait_0 & ((ramiframload_1))) # (!ccifiwait_0 & (instr[1]))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(instr[1]),
	.datad(ramiframload_1),
	.cin(gnd),
	.combout(dcifimemload_1),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[1]~21 .lut_mask = 16'hFA50;
defparam \dcif.imemload[1]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N24
cycloneive_lcell_comb \dcif.imemload[15]~22 (
// Equation(s):
// dcifimemload_15 = (ccifiwait_0 & (ramiframload_15)) # (!ccifiwait_0 & ((instr[15])))

	.dataa(gnd),
	.datab(ramiframload_15),
	.datac(instr[15]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_15),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[15]~22 .lut_mask = 16'hCCF0;
defparam \dcif.imemload[15]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N4
cycloneive_lcell_comb \dcif.imemload[14]~23 (
// Equation(s):
// dcifimemload_14 = (ccifiwait_0 & (ramiframload_14)) # (!ccifiwait_0 & ((instr[14])))

	.dataa(ccifiwait_0),
	.datab(ramiframload_14),
	.datac(instr[14]),
	.datad(gnd),
	.cin(gnd),
	.combout(dcifimemload_14),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[14]~23 .lut_mask = 16'hD8D8;
defparam \dcif.imemload[14]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N14
cycloneive_lcell_comb \dcif.imemload[13]~24 (
// Equation(s):
// dcifimemload_13 = (ccifiwait_0 & ((ramiframload_13))) # (!ccifiwait_0 & (instr[13]))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[13]),
	.datad(ramiframload_13),
	.cin(gnd),
	.combout(dcifimemload_13),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[13]~24 .lut_mask = 16'hFC30;
defparam \dcif.imemload[13]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N14
cycloneive_lcell_comb \dcif.imemload[12]~25 (
// Equation(s):
// dcifimemload_12 = (ccifiwait_0 & ((ramiframload_12))) # (!ccifiwait_0 & (instr[12]))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(instr[12]),
	.datad(ramiframload_12),
	.cin(gnd),
	.combout(dcifimemload_12),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[12]~25 .lut_mask = 16'hFA50;
defparam \dcif.imemload[12]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N20
cycloneive_lcell_comb \dcif.imemload[11]~26 (
// Equation(s):
// dcifimemload_11 = (ccifiwait_0 & ((ramiframload_11))) # (!ccifiwait_0 & (instr[11]))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[11]),
	.datad(ramiframload_11),
	.cin(gnd),
	.combout(dcifimemload_11),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[11]~26 .lut_mask = 16'hFC30;
defparam \dcif.imemload[11]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N0
cycloneive_lcell_comb \dcif.imemload[10]~27 (
// Equation(s):
// dcifimemload_10 = (ccifiwait_0 & (ramiframload_10)) # (!ccifiwait_0 & ((instr[10])))

	.dataa(ramiframload_10),
	.datab(gnd),
	.datac(instr[10]),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(dcifimemload_10),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[10]~27 .lut_mask = 16'hAAF0;
defparam \dcif.imemload[10]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N14
cycloneive_lcell_comb \dcif.imemload[9]~28 (
// Equation(s):
// dcifimemload_9 = (ccifiwait_0 & ((ramiframload_9))) # (!ccifiwait_0 & (instr[9]))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[9]),
	.datad(ramiframload_9),
	.cin(gnd),
	.combout(dcifimemload_9),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[9]~28 .lut_mask = 16'hFC30;
defparam \dcif.imemload[9]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N24
cycloneive_lcell_comb \dcif.imemload[8]~29 (
// Equation(s):
// dcifimemload_8 = (ccifiwait_0 & ((ramiframload_8))) # (!ccifiwait_0 & (instr[8]))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[8]),
	.datad(ramiframload_8),
	.cin(gnd),
	.combout(dcifimemload_8),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[8]~29 .lut_mask = 16'hFC30;
defparam \dcif.imemload[8]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N16
cycloneive_lcell_comb \dcif.imemload[7]~30 (
// Equation(s):
// dcifimemload_7 = (ccifiwait_0 & ((ramiframload_7))) # (!ccifiwait_0 & (instr[7]))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(instr[7]),
	.datad(ramiframload_7),
	.cin(gnd),
	.combout(dcifimemload_7),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[7]~30 .lut_mask = 16'hFA50;
defparam \dcif.imemload[7]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N22
cycloneive_lcell_comb \dcif.imemload[6]~31 (
// Equation(s):
// dcifimemload_6 = (ccifiwait_0 & ((ramiframload_6))) # (!ccifiwait_0 & (instr[6]))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(instr[6]),
	.datad(ramiframload_6),
	.cin(gnd),
	.combout(dcifimemload_6),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[6]~31 .lut_mask = 16'hFC30;
defparam \dcif.imemload[6]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N18
cycloneive_lcell_comb \dcif.dhit~0 (
// Equation(s):
// dcifdhit = (always1 & ((reg_WEN1) # (reg_REN1)))

	.dataa(gnd),
	.datab(always1),
	.datac(reg_WEN),
	.datad(reg_REN),
	.cin(gnd),
	.combout(dcifdhit),
	.cout());
// synopsys translate_off
defparam \dcif.dhit~0 .lut_mask = 16'hCCC0;
defparam \dcif.dhit~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N24
cycloneive_lcell_comb \daddr~0 (
// Equation(s):
// \daddr~0_combout  = (\nRST~input_o  & Selector30)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Selector30),
	.cin(gnd),
	.combout(\daddr~0_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~0 .lut_mask = 16'hF000;
defparam \daddr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N20
cycloneive_lcell_comb \daddr[1]~1 (
// Equation(s):
// \daddr[1]~1_combout  = ((!reg_REN1 & (!reg_WEN1 & always1))) # (!\nRST~input_o )

	.dataa(nRST),
	.datab(reg_REN),
	.datac(reg_WEN),
	.datad(always1),
	.cin(gnd),
	.combout(\daddr[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \daddr[1]~1 .lut_mask = 16'h5755;
defparam \daddr[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N26
cycloneive_lcell_comb \daddr~2 (
// Equation(s):
// \daddr~2_combout  = (\nRST~input_o  & ((Selector31) # ((ShiftRight0 & Selector24))))

	.dataa(ShiftRight0),
	.datab(Selector31),
	.datac(nRST),
	.datad(Selector24),
	.cin(gnd),
	.combout(\daddr~2_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~2 .lut_mask = 16'hE0C0;
defparam \daddr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N12
cycloneive_lcell_comb \daddr~3 (
// Equation(s):
// \daddr~3_combout  = (\nRST~input_o  & Selector28)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Selector28),
	.cin(gnd),
	.combout(\daddr~3_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~3 .lut_mask = 16'hF000;
defparam \daddr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N30
cycloneive_lcell_comb \daddr~4 (
// Equation(s):
// \daddr~4_combout  = (\nRST~input_o  & ((Selector29) # ((ShiftRight03 & Selector22))))

	.dataa(ShiftRight03),
	.datab(Selector22),
	.datac(nRST),
	.datad(Selector29),
	.cin(gnd),
	.combout(\daddr~4_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~4 .lut_mask = 16'hF080;
defparam \daddr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N22
cycloneive_lcell_comb \daddr~5 (
// Equation(s):
// \daddr~5_combout  = (\nRST~input_o  & ((Selector26) # ((Selector241 & ShiftLeft0))))

	.dataa(Selector26),
	.datab(Selector241),
	.datac(ShiftLeft0),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~5_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~5 .lut_mask = 16'hEA00;
defparam \daddr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N0
cycloneive_lcell_comb \daddr~6 (
// Equation(s):
// \daddr~6_combout  = (\nRST~input_o  & Selector27)

	.dataa(nRST),
	.datab(gnd),
	.datac(gnd),
	.datad(Selector27),
	.cin(gnd),
	.combout(\daddr~6_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~6 .lut_mask = 16'hAA00;
defparam \daddr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N4
cycloneive_lcell_comb \daddr~7 (
// Equation(s):
// \daddr~7_combout  = (Selector242 & \nRST~input_o )

	.dataa(gnd),
	.datab(Selector242),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~7_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~7 .lut_mask = 16'hCC00;
defparam \daddr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N26
cycloneive_lcell_comb \daddr~8 (
// Equation(s):
// \daddr~8_combout  = (\nRST~input_o  & Selector25)

	.dataa(gnd),
	.datab(nRST),
	.datac(Selector25),
	.datad(gnd),
	.cin(gnd),
	.combout(\daddr~8_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~8 .lut_mask = 16'hC0C0;
defparam \daddr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N28
cycloneive_lcell_comb \daddr~9 (
// Equation(s):
// \daddr~9_combout  = (\nRST~input_o  & Selector221)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(Selector221),
	.cin(gnd),
	.combout(\daddr~9_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~9 .lut_mask = 16'hCC00;
defparam \daddr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N14
cycloneive_lcell_comb \daddr~10 (
// Equation(s):
// \daddr~10_combout  = (\nRST~input_o  & ((Selector232) # ((Selector23) # (Selector231))))

	.dataa(nRST),
	.datab(Selector232),
	.datac(Selector23),
	.datad(Selector231),
	.cin(gnd),
	.combout(\daddr~10_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~10 .lut_mask = 16'hAAA8;
defparam \daddr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N12
cycloneive_lcell_comb \daddr~11 (
// Equation(s):
// \daddr~11_combout  = (\nRST~input_o  & ((Selector201) # ((Selector202) # (Selector20))))

	.dataa(nRST),
	.datab(Selector201),
	.datac(Selector202),
	.datad(Selector20),
	.cin(gnd),
	.combout(\daddr~11_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~11 .lut_mask = 16'hAAA8;
defparam \daddr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N24
cycloneive_lcell_comb \daddr~12 (
// Equation(s):
// \daddr~12_combout  = (\nRST~input_o  & ((Selector21) # ((Selector212) # (Selector211))))

	.dataa(Selector21),
	.datab(nRST),
	.datac(Selector212),
	.datad(Selector211),
	.cin(gnd),
	.combout(\daddr~12_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~12 .lut_mask = 16'hCCC8;
defparam \daddr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N20
cycloneive_lcell_comb \daddr~13 (
// Equation(s):
// \daddr~13_combout  = (Selector18 & \nRST~input_o )

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector18),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~13_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~13 .lut_mask = 16'hF000;
defparam \daddr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N14
cycloneive_lcell_comb \daddr~14 (
// Equation(s):
// \daddr~14_combout  = (Selector19 & \nRST~input_o )

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector19),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~14_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~14 .lut_mask = 16'hF000;
defparam \daddr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N28
cycloneive_lcell_comb \daddr~15 (
// Equation(s):
// \daddr~15_combout  = (\nRST~input_o  & Selector16)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Selector16),
	.cin(gnd),
	.combout(\daddr~15_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~15 .lut_mask = 16'hF000;
defparam \daddr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N30
cycloneive_lcell_comb \daddr~16 (
// Equation(s):
// \daddr~16_combout  = (\nRST~input_o  & Selector17)

	.dataa(gnd),
	.datab(nRST),
	.datac(Selector17),
	.datad(gnd),
	.cin(gnd),
	.combout(\daddr~16_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~16 .lut_mask = 16'hC0C0;
defparam \daddr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N2
cycloneive_lcell_comb \daddr~17 (
// Equation(s):
// \daddr~17_combout  = (\nRST~input_o  & ((Selector14) # ((Selector141) # (Selector142))))

	.dataa(nRST),
	.datab(Selector14),
	.datac(Selector141),
	.datad(Selector142),
	.cin(gnd),
	.combout(\daddr~17_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~17 .lut_mask = 16'hAAA8;
defparam \daddr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N4
cycloneive_lcell_comb \daddr~18 (
// Equation(s):
// \daddr~18_combout  = (\nRST~input_o  & Selector15)

	.dataa(nRST),
	.datab(gnd),
	.datac(gnd),
	.datad(Selector15),
	.cin(gnd),
	.combout(\daddr~18_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~18 .lut_mask = 16'hAA00;
defparam \daddr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N16
cycloneive_lcell_comb \daddr~19 (
// Equation(s):
// \daddr~19_combout  = (Selector12 & \nRST~input_o )

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector12),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~19_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~19 .lut_mask = 16'hF000;
defparam \daddr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N24
cycloneive_lcell_comb \daddr~20 (
// Equation(s):
// \daddr~20_combout  = (Selector13 & \nRST~input_o )

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector13),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~20_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~20 .lut_mask = 16'hF000;
defparam \daddr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N4
cycloneive_lcell_comb \daddr~21 (
// Equation(s):
// \daddr~21_combout  = (\nRST~input_o  & ((Selector101) # ((Selector10) # (Selector102))))

	.dataa(nRST),
	.datab(Selector101),
	.datac(Selector10),
	.datad(Selector102),
	.cin(gnd),
	.combout(\daddr~21_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~21 .lut_mask = 16'hAAA8;
defparam \daddr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N30
cycloneive_lcell_comb \daddr~22 (
// Equation(s):
// \daddr~22_combout  = (\nRST~input_o  & ((Selector11) # ((ShiftRight01 & Selector8))))

	.dataa(Selector11),
	.datab(nRST),
	.datac(ShiftRight01),
	.datad(Selector8),
	.cin(gnd),
	.combout(\daddr~22_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~22 .lut_mask = 16'hC888;
defparam \daddr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N14
cycloneive_lcell_comb \daddr~23 (
// Equation(s):
// \daddr~23_combout  = (\nRST~input_o  & ((Selector81) # ((Selector83) # (Selector82))))

	.dataa(nRST),
	.datab(Selector81),
	.datac(Selector83),
	.datad(Selector82),
	.cin(gnd),
	.combout(\daddr~23_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~23 .lut_mask = 16'hAAA8;
defparam \daddr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N4
cycloneive_lcell_comb \daddr~24 (
// Equation(s):
// \daddr~24_combout  = (\nRST~input_o  & ((Selector91) # ((Selector9) # (Selector92))))

	.dataa(nRST),
	.datab(Selector91),
	.datac(Selector9),
	.datad(Selector92),
	.cin(gnd),
	.combout(\daddr~24_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~24 .lut_mask = 16'hAAA8;
defparam \daddr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N4
cycloneive_lcell_comb \daddr~25 (
// Equation(s):
// \daddr~25_combout  = (\nRST~input_o  & Selector6)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(Selector6),
	.cin(gnd),
	.combout(\daddr~25_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~25 .lut_mask = 16'hCC00;
defparam \daddr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N26
cycloneive_lcell_comb \daddr~26 (
// Equation(s):
// \daddr~26_combout  = (Selector7 & \nRST~input_o )

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector7),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~26_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~26 .lut_mask = 16'hF000;
defparam \daddr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N28
cycloneive_lcell_comb \daddr~27 (
// Equation(s):
// \daddr~27_combout  = (\nRST~input_o  & Selector41)

	.dataa(gnd),
	.datab(nRST),
	.datac(Selector41),
	.datad(gnd),
	.cin(gnd),
	.combout(\daddr~27_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~27 .lut_mask = 16'hC0C0;
defparam \daddr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N4
cycloneive_lcell_comb \daddr~28 (
// Equation(s):
// \daddr~28_combout  = (\nRST~input_o  & ((Selector5) # ((Selector4 & ShiftRight02))))

	.dataa(Selector4),
	.datab(ShiftRight02),
	.datac(Selector5),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~28_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~28 .lut_mask = 16'hF800;
defparam \daddr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N24
cycloneive_lcell_comb \daddr~29 (
// Equation(s):
// \daddr~29_combout  = (\nRST~input_o  & Selector2)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Selector2),
	.cin(gnd),
	.combout(\daddr~29_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~29 .lut_mask = 16'hF000;
defparam \daddr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N12
cycloneive_lcell_comb \daddr~30 (
// Equation(s):
// \daddr~30_combout  = (\nRST~input_o  & Selector3)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(Selector3),
	.cin(gnd),
	.combout(\daddr~30_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~30 .lut_mask = 16'hCC00;
defparam \daddr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N16
cycloneive_lcell_comb \daddr~31 (
// Equation(s):
// \daddr~31_combout  = (\nRST~input_o  & Selector0)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(Selector0),
	.cin(gnd),
	.combout(\daddr~31_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~31 .lut_mask = 16'hCC00;
defparam \daddr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N8
cycloneive_lcell_comb \daddr~32 (
// Equation(s):
// \daddr~32_combout  = (\nRST~input_o  & Selector1)

	.dataa(nRST),
	.datab(gnd),
	.datac(Selector1),
	.datad(gnd),
	.cin(gnd),
	.combout(\daddr~32_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~32 .lut_mask = 16'hA0A0;
defparam \daddr~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N22
cycloneive_lcell_comb \instr~0 (
// Equation(s):
// \instr~0_combout  = (\nRST~input_o  & ramiframload_30)

	.dataa(nRST),
	.datab(ramiframload_30),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr~0_combout ),
	.cout());
// synopsys translate_off
defparam \instr~0 .lut_mask = 16'h8888;
defparam \instr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N4
cycloneive_lcell_comb \instr~1 (
// Equation(s):
// \instr~1_combout  = (ramiframload_31 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_31),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~1_combout ),
	.cout());
// synopsys translate_off
defparam \instr~1 .lut_mask = 16'hCC00;
defparam \instr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N12
cycloneive_lcell_comb \instr~2 (
// Equation(s):
// \instr~2_combout  = (ramiframload_27 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_27),
	.datac(nRST),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr~2_combout ),
	.cout());
// synopsys translate_off
defparam \instr~2 .lut_mask = 16'hC0C0;
defparam \instr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N8
cycloneive_lcell_comb \instr~3 (
// Equation(s):
// \instr~3_combout  = (ramiframload_26 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_26),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~3_combout ),
	.cout());
// synopsys translate_off
defparam \instr~3 .lut_mask = 16'hCC00;
defparam \instr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N30
cycloneive_lcell_comb \instr~4 (
// Equation(s):
// \instr~4_combout  = (\nRST~input_o  & ramiframload_29)

	.dataa(nRST),
	.datab(gnd),
	.datac(ramiframload_29),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr~4_combout ),
	.cout());
// synopsys translate_off
defparam \instr~4 .lut_mask = 16'hA0A0;
defparam \instr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N6
cycloneive_lcell_comb \instr~5 (
// Equation(s):
// \instr~5_combout  = (\nRST~input_o  & ramiframload_28)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(ramiframload_28),
	.cin(gnd),
	.combout(\instr~5_combout ),
	.cout());
// synopsys translate_off
defparam \instr~5 .lut_mask = 16'hCC00;
defparam \instr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N10
cycloneive_lcell_comb \instr~6 (
// Equation(s):
// \instr~6_combout  = (\nRST~input_o  & ramiframload_19)

	.dataa(nRST),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_19),
	.cin(gnd),
	.combout(\instr~6_combout ),
	.cout());
// synopsys translate_off
defparam \instr~6 .lut_mask = 16'hAA00;
defparam \instr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N21
dffeas \instr[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[19]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[19] .is_wysiwyg = "true";
defparam \instr[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N30
cycloneive_lcell_comb \instr~7 (
// Equation(s):
// \instr~7_combout  = (\nRST~input_o  & ramiframload_18)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(ramiframload_18),
	.cin(gnd),
	.combout(\instr~7_combout ),
	.cout());
// synopsys translate_off
defparam \instr~7 .lut_mask = 16'hCC00;
defparam \instr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N29
dffeas \instr[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~7_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[18]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[18] .is_wysiwyg = "true";
defparam \instr[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N16
cycloneive_lcell_comb \instr~8 (
// Equation(s):
// \instr~8_combout  = (\nRST~input_o  & ramiframload_16)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(ramiframload_16),
	.cin(gnd),
	.combout(\instr~8_combout ),
	.cout());
// synopsys translate_off
defparam \instr~8 .lut_mask = 16'hCC00;
defparam \instr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N24
cycloneive_lcell_comb \instr[16]~feeder (
// Equation(s):
// \instr[16]~feeder_combout  = \instr~8_combout 

	.dataa(gnd),
	.datab(\instr~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[16]~feeder .lut_mask = 16'hCCCC;
defparam \instr[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N16
cycloneive_lcell_comb \instr~9 (
// Equation(s):
// \instr~9_combout  = (ramiframload_17 & \nRST~input_o )

	.dataa(ramiframload_17),
	.datab(nRST),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr~9_combout ),
	.cout());
// synopsys translate_off
defparam \instr~9 .lut_mask = 16'h8888;
defparam \instr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N4
cycloneive_lcell_comb \instr~10 (
// Equation(s):
// \instr~10_combout  = (ramiframload_20 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_20),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~10_combout ),
	.cout());
// synopsys translate_off
defparam \instr~10 .lut_mask = 16'hCC00;
defparam \instr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N19
dffeas \instr[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[20]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[20] .is_wysiwyg = "true";
defparam \instr[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N20
cycloneive_lcell_comb \instr~11 (
// Equation(s):
// \instr~11_combout  = (\nRST~input_o  & ramiframload_24)

	.dataa(gnd),
	.datab(nRST),
	.datac(ramiframload_24),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr~11_combout ),
	.cout());
// synopsys translate_off
defparam \instr~11 .lut_mask = 16'hC0C0;
defparam \instr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N15
dffeas \instr[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[24]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[24] .is_wysiwyg = "true";
defparam \instr[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N6
cycloneive_lcell_comb \instr~12 (
// Equation(s):
// \instr~12_combout  = (ramiframload_23 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_23),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~12_combout ),
	.cout());
// synopsys translate_off
defparam \instr~12 .lut_mask = 16'hCC00;
defparam \instr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N1
dffeas \instr[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~12_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[23]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[23] .is_wysiwyg = "true";
defparam \instr[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N24
cycloneive_lcell_comb \instr~13 (
// Equation(s):
// \instr~13_combout  = (\nRST~input_o  & ramiframload_21)

	.dataa(nRST),
	.datab(gnd),
	.datac(ramiframload_21),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr~13_combout ),
	.cout());
// synopsys translate_off
defparam \instr~13 .lut_mask = 16'hA0A0;
defparam \instr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y37_N1
dffeas \instr[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~13_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[21]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[21] .is_wysiwyg = "true";
defparam \instr[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N22
cycloneive_lcell_comb \instr~14 (
// Equation(s):
// \instr~14_combout  = (\nRST~input_o  & ramiframload_22)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(ramiframload_22),
	.cin(gnd),
	.combout(\instr~14_combout ),
	.cout());
// synopsys translate_off
defparam \instr~14 .lut_mask = 16'hCC00;
defparam \instr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N17
dffeas \instr[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~14_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[22]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[22] .is_wysiwyg = "true";
defparam \instr[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N18
cycloneive_lcell_comb \instr~15 (
// Equation(s):
// \instr~15_combout  = (\nRST~input_o  & ramiframload_25)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(ramiframload_25),
	.cin(gnd),
	.combout(\instr~15_combout ),
	.cout());
// synopsys translate_off
defparam \instr~15 .lut_mask = 16'hF000;
defparam \instr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N11
dffeas \instr[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~15_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[25]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[25] .is_wysiwyg = "true";
defparam \instr[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N4
cycloneive_lcell_comb \instr~16 (
// Equation(s):
// \instr~16_combout  = (ramiframload_3 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_3),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~16_combout ),
	.cout());
// synopsys translate_off
defparam \instr~16 .lut_mask = 16'hCC00;
defparam \instr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y29_N1
dffeas \instr[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~16_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[3]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[3] .is_wysiwyg = "true";
defparam \instr[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N10
cycloneive_lcell_comb \instr~17 (
// Equation(s):
// \instr~17_combout  = (\nRST~input_o  & ramiframload_4)

	.dataa(nRST),
	.datab(gnd),
	.datac(ramiframload_4),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr~17_combout ),
	.cout());
// synopsys translate_off
defparam \instr~17 .lut_mask = 16'hA0A0;
defparam \instr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N25
dffeas \instr[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~17_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[4]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[4] .is_wysiwyg = "true";
defparam \instr[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N28
cycloneive_lcell_comb \instr~18 (
// Equation(s):
// \instr~18_combout  = (ramiframload_2 & \nRST~input_o )

	.dataa(gnd),
	.datab(gnd),
	.datac(ramiframload_2),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~18_combout ),
	.cout());
// synopsys translate_off
defparam \instr~18 .lut_mask = 16'hF000;
defparam \instr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y29_N31
dffeas \instr[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~18_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[2]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[2] .is_wysiwyg = "true";
defparam \instr[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N26
cycloneive_lcell_comb \instr~19 (
// Equation(s):
// \instr~19_combout  = (ramiframload_5 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_5),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~19_combout ),
	.cout());
// synopsys translate_off
defparam \instr~19 .lut_mask = 16'hCC00;
defparam \instr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N17
dffeas \instr[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~19_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[5]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[5] .is_wysiwyg = "true";
defparam \instr[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N28
cycloneive_lcell_comb \instr~20 (
// Equation(s):
// \instr~20_combout  = (\nRST~input_o  & ramiframload_0)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(ramiframload_0),
	.cin(gnd),
	.combout(\instr~20_combout ),
	.cout());
// synopsys translate_off
defparam \instr~20 .lut_mask = 16'hCC00;
defparam \instr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y30_N31
dffeas \instr[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~20_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[0]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[0] .is_wysiwyg = "true";
defparam \instr[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N2
cycloneive_lcell_comb \instr~21 (
// Equation(s):
// \instr~21_combout  = (\nRST~input_o  & ramiframload_1)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(ramiframload_1),
	.cin(gnd),
	.combout(\instr~21_combout ),
	.cout());
// synopsys translate_off
defparam \instr~21 .lut_mask = 16'hCC00;
defparam \instr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y30_N29
dffeas \instr[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~21_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[1]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[1] .is_wysiwyg = "true";
defparam \instr[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N28
cycloneive_lcell_comb \instr~22 (
// Equation(s):
// \instr~22_combout  = (ramiframload_15 & \nRST~input_o )

	.dataa(gnd),
	.datab(gnd),
	.datac(ramiframload_15),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~22_combout ),
	.cout());
// synopsys translate_off
defparam \instr~22 .lut_mask = 16'hF000;
defparam \instr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N25
dffeas \instr[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~22_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[15]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[15] .is_wysiwyg = "true";
defparam \instr[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N26
cycloneive_lcell_comb \instr~23 (
// Equation(s):
// \instr~23_combout  = (\nRST~input_o  & ramiframload_14)

	.dataa(nRST),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_14),
	.cin(gnd),
	.combout(\instr~23_combout ),
	.cout());
// synopsys translate_off
defparam \instr~23 .lut_mask = 16'hAA00;
defparam \instr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N5
dffeas \instr[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~23_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[14]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[14] .is_wysiwyg = "true";
defparam \instr[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N16
cycloneive_lcell_comb \instr~24 (
// Equation(s):
// \instr~24_combout  = (\nRST~input_o  & ramiframload_13)

	.dataa(nRST),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_13),
	.cin(gnd),
	.combout(\instr~24_combout ),
	.cout());
// synopsys translate_off
defparam \instr~24 .lut_mask = 16'hAA00;
defparam \instr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N15
dffeas \instr[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~24_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[13]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[13] .is_wysiwyg = "true";
defparam \instr[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N2
cycloneive_lcell_comb \instr~25 (
// Equation(s):
// \instr~25_combout  = (ramiframload_12 & \nRST~input_o )

	.dataa(ramiframload_12),
	.datab(gnd),
	.datac(nRST),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr~25_combout ),
	.cout());
// synopsys translate_off
defparam \instr~25 .lut_mask = 16'hA0A0;
defparam \instr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N15
dffeas \instr[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[12]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[12] .is_wysiwyg = "true";
defparam \instr[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N26
cycloneive_lcell_comb \instr~26 (
// Equation(s):
// \instr~26_combout  = (\nRST~input_o  & ramiframload_11)

	.dataa(nRST),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_11),
	.cin(gnd),
	.combout(\instr~26_combout ),
	.cout());
// synopsys translate_off
defparam \instr~26 .lut_mask = 16'hAA00;
defparam \instr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N21
dffeas \instr[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~26_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[11]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[11] .is_wysiwyg = "true";
defparam \instr[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N12
cycloneive_lcell_comb \instr~27 (
// Equation(s):
// \instr~27_combout  = (ramiframload_10 & \nRST~input_o )

	.dataa(gnd),
	.datab(gnd),
	.datac(ramiframload_10),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~27_combout ),
	.cout());
// synopsys translate_off
defparam \instr~27 .lut_mask = 16'hF000;
defparam \instr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N1
dffeas \instr[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~27_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[10]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[10] .is_wysiwyg = "true";
defparam \instr[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N6
cycloneive_lcell_comb \instr~28 (
// Equation(s):
// \instr~28_combout  = (\nRST~input_o  & ramiframload_9)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(ramiframload_9),
	.cin(gnd),
	.combout(\instr~28_combout ),
	.cout());
// synopsys translate_off
defparam \instr~28 .lut_mask = 16'hCC00;
defparam \instr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N15
dffeas \instr[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~28_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[9]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[9] .is_wysiwyg = "true";
defparam \instr[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N14
cycloneive_lcell_comb \instr~29 (
// Equation(s):
// \instr~29_combout  = (\nRST~input_o  & ramiframload_8)

	.dataa(nRST),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_8),
	.cin(gnd),
	.combout(\instr~29_combout ),
	.cout());
// synopsys translate_off
defparam \instr~29 .lut_mask = 16'hAA00;
defparam \instr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N25
dffeas \instr[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~29_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[8]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[8] .is_wysiwyg = "true";
defparam \instr[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N8
cycloneive_lcell_comb \instr~30 (
// Equation(s):
// \instr~30_combout  = (\nRST~input_o  & ramiframload_7)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(ramiframload_7),
	.cin(gnd),
	.combout(\instr~30_combout ),
	.cout());
// synopsys translate_off
defparam \instr~30 .lut_mask = 16'hF000;
defparam \instr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N17
dffeas \instr[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~30_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[7]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[7] .is_wysiwyg = "true";
defparam \instr[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N6
cycloneive_lcell_comb \instr~31 (
// Equation(s):
// \instr~31_combout  = (ramiframload_6 & \nRST~input_o )

	.dataa(gnd),
	.datab(ramiframload_6),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~31_combout ),
	.cout());
// synopsys translate_off
defparam \instr~31 .lut_mask = 16'hCC00;
defparam \instr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N23
dffeas \instr[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~31_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[6]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[6] .is_wysiwyg = "true";
defparam \instr[6] .power_up = "low";
// synopsys translate_on

endmodule

module datapath (
	PC_29,
	PC_28,
	PC_31,
	PC_30,
	dpifhalt,
	PC_1,
	reg_WEN,
	reg_REN,
	PC_0,
	PC_3,
	PC_2,
	PC_5,
	PC_4,
	PC_7,
	PC_6,
	PC_9,
	PC_8,
	PC_11,
	PC_10,
	PC_13,
	PC_12,
	PC_15,
	PC_14,
	PC_17,
	PC_16,
	PC_19,
	PC_18,
	PC_21,
	PC_20,
	PC_23,
	PC_22,
	PC_25,
	PC_24,
	PC_27,
	PC_26,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	instr_30,
	ccifiwait_0,
	dcifimemload_30,
	instr_31,
	dcifimemload_31,
	instr_27,
	dcifimemload_27,
	instr_26,
	dcifimemload_26,
	instr_29,
	dcifimemload_29,
	instr_28,
	dcifimemload_28,
	dcifimemload_19,
	dcifimemload_18,
	instr_16,
	dcifimemload_16,
	instr_17,
	dcifimemload_17,
	Mux63,
	Mux631,
	dcifimemload_20,
	dcifimemload_24,
	dcifimemload_23,
	dcifimemload_21,
	dcifimemload_22,
	dcifimemload_25,
	dcifimemload_3,
	dcifimemload_4,
	dcifimemload_2,
	dcifimemload_5,
	dcifimemload_0,
	dcifimemload_1,
	dcifimemload_15,
	Mux32,
	Mux321,
	Mux33,
	Mux331,
	Mux34,
	Mux341,
	Mux35,
	Mux351,
	Mux36,
	Mux361,
	Mux37,
	Mux371,
	Mux38,
	Mux381,
	Mux39,
	Mux391,
	Mux40,
	Mux401,
	Mux41,
	Mux411,
	Mux42,
	Mux421,
	Mux43,
	Mux431,
	Mux44,
	Mux441,
	Mux45,
	Mux451,
	Mux46,
	Mux461,
	Mux47,
	Mux471,
	Mux48,
	Mux481,
	dcifimemload_14,
	Mux49,
	Mux491,
	dcifimemload_13,
	Mux50,
	Mux501,
	dcifimemload_12,
	Mux51,
	Mux511,
	dcifimemload_11,
	Mux52,
	Mux521,
	dcifimemload_10,
	Mux53,
	Mux531,
	dcifimemload_9,
	Mux54,
	Mux541,
	dcifimemload_8,
	Mux55,
	Mux551,
	dcifimemload_7,
	Mux56,
	Mux561,
	dcifimemload_6,
	Mux57,
	Mux571,
	Mux58,
	Mux581,
	Mux59,
	Mux591,
	Mux60,
	Mux601,
	Mux61,
	Mux611,
	Mux62,
	Mux621,
	Selector31,
	ShiftRight0,
	Selector24,
	Selector8,
	Selector0,
	Selector3,
	Selector4,
	Selector7,
	Selector11,
	ShiftRight01,
	Selector15,
	Selector22,
	Selector28,
	Selector29,
	ShiftRight02,
	ShiftRight03,
	ShiftLeft0,
	Selector10,
	Selector101,
	Selector102,
	Selector2,
	Selector1,
	Selector41,
	Selector5,
	Selector12,
	Selector241,
	Selector242,
	Selector13,
	Selector25,
	Selector14,
	Selector141,
	Selector142,
	Selector27,
	Selector16,
	Selector18,
	Selector17,
	Selector6,
	Selector26,
	Selector19,
	Selector20,
	Selector201,
	Selector202,
	Selector21,
	Selector211,
	Selector212,
	Selector81,
	Selector82,
	Selector83,
	Selector9,
	Selector91,
	Selector92,
	Selector221,
	Selector30,
	Selector23,
	Selector231,
	Selector232,
	dcifdhit,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
output 	PC_29;
output 	PC_28;
output 	PC_31;
output 	PC_30;
output 	dpifhalt;
output 	PC_1;
output 	reg_WEN;
output 	reg_REN;
output 	PC_0;
output 	PC_3;
output 	PC_2;
output 	PC_5;
output 	PC_4;
output 	PC_7;
output 	PC_6;
output 	PC_9;
output 	PC_8;
output 	PC_11;
output 	PC_10;
output 	PC_13;
output 	PC_12;
output 	PC_15;
output 	PC_14;
output 	PC_17;
output 	PC_16;
output 	PC_19;
output 	PC_18;
output 	PC_21;
output 	PC_20;
output 	PC_23;
output 	PC_22;
output 	PC_25;
output 	PC_24;
output 	PC_27;
output 	PC_26;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	instr_30;
input 	ccifiwait_0;
input 	dcifimemload_30;
input 	instr_31;
input 	dcifimemload_31;
input 	instr_27;
input 	dcifimemload_27;
input 	instr_26;
input 	dcifimemload_26;
input 	instr_29;
input 	dcifimemload_29;
input 	instr_28;
input 	dcifimemload_28;
input 	dcifimemload_19;
input 	dcifimemload_18;
input 	instr_16;
input 	dcifimemload_16;
input 	instr_17;
input 	dcifimemload_17;
output 	Mux63;
output 	Mux631;
input 	dcifimemload_20;
input 	dcifimemload_24;
input 	dcifimemload_23;
input 	dcifimemload_21;
input 	dcifimemload_22;
input 	dcifimemload_25;
input 	dcifimemload_3;
input 	dcifimemload_4;
input 	dcifimemload_2;
input 	dcifimemload_5;
input 	dcifimemload_0;
input 	dcifimemload_1;
input 	dcifimemload_15;
output 	Mux32;
output 	Mux321;
output 	Mux33;
output 	Mux331;
output 	Mux34;
output 	Mux341;
output 	Mux35;
output 	Mux351;
output 	Mux36;
output 	Mux361;
output 	Mux37;
output 	Mux371;
output 	Mux38;
output 	Mux381;
output 	Mux39;
output 	Mux391;
output 	Mux40;
output 	Mux401;
output 	Mux41;
output 	Mux411;
output 	Mux42;
output 	Mux421;
output 	Mux43;
output 	Mux431;
output 	Mux44;
output 	Mux441;
output 	Mux45;
output 	Mux451;
output 	Mux46;
output 	Mux461;
output 	Mux47;
output 	Mux471;
output 	Mux48;
output 	Mux481;
input 	dcifimemload_14;
output 	Mux49;
output 	Mux491;
input 	dcifimemload_13;
output 	Mux50;
output 	Mux501;
input 	dcifimemload_12;
output 	Mux51;
output 	Mux511;
input 	dcifimemload_11;
output 	Mux52;
output 	Mux521;
input 	dcifimemload_10;
output 	Mux53;
output 	Mux531;
input 	dcifimemload_9;
output 	Mux54;
output 	Mux541;
input 	dcifimemload_8;
output 	Mux55;
output 	Mux551;
input 	dcifimemload_7;
output 	Mux56;
output 	Mux561;
input 	dcifimemload_6;
output 	Mux57;
output 	Mux571;
output 	Mux58;
output 	Mux581;
output 	Mux59;
output 	Mux591;
output 	Mux60;
output 	Mux601;
output 	Mux61;
output 	Mux611;
output 	Mux62;
output 	Mux621;
output 	Selector31;
output 	ShiftRight0;
output 	Selector24;
output 	Selector8;
output 	Selector0;
output 	Selector3;
output 	Selector4;
output 	Selector7;
output 	Selector11;
output 	ShiftRight01;
output 	Selector15;
output 	Selector22;
output 	Selector28;
output 	Selector29;
output 	ShiftRight02;
output 	ShiftRight03;
output 	ShiftLeft0;
output 	Selector10;
output 	Selector101;
output 	Selector102;
output 	Selector2;
output 	Selector1;
output 	Selector41;
output 	Selector5;
output 	Selector12;
output 	Selector241;
output 	Selector242;
output 	Selector13;
output 	Selector25;
output 	Selector14;
output 	Selector141;
output 	Selector142;
output 	Selector27;
output 	Selector16;
output 	Selector18;
output 	Selector17;
output 	Selector6;
output 	Selector26;
output 	Selector19;
output 	Selector20;
output 	Selector201;
output 	Selector202;
output 	Selector21;
output 	Selector211;
output 	Selector212;
output 	Selector81;
output 	Selector82;
output 	Selector83;
output 	Selector9;
output 	Selector91;
output 	Selector92;
output 	Selector221;
output 	Selector30;
output 	Selector23;
output 	Selector231;
output 	Selector232;
input 	dcifdhit;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add0~1 ;
wire \Add0~0_combout ;
wire \Add0~3 ;
wire \Add0~2_combout ;
wire \Add0~5 ;
wire \Add0~4_combout ;
wire \Add0~7 ;
wire \Add0~6_combout ;
wire \Add0~9 ;
wire \Add0~8_combout ;
wire \Add0~11 ;
wire \Add0~10_combout ;
wire \Add0~13 ;
wire \Add0~12_combout ;
wire \Add0~15 ;
wire \Add0~14_combout ;
wire \Add0~17 ;
wire \Add0~16_combout ;
wire \Add0~19 ;
wire \Add0~18_combout ;
wire \Add0~21 ;
wire \Add0~20_combout ;
wire \Add0~23 ;
wire \Add0~22_combout ;
wire \Add0~25 ;
wire \Add0~24_combout ;
wire \Add0~27 ;
wire \Add0~26_combout ;
wire \Add0~29 ;
wire \Add0~28_combout ;
wire \Add0~31 ;
wire \Add0~30_combout ;
wire \Add0~33 ;
wire \Add0~32_combout ;
wire \Add0~35 ;
wire \Add0~34_combout ;
wire \Add0~37 ;
wire \Add0~36_combout ;
wire \Add0~39 ;
wire \Add0~38_combout ;
wire \Add0~41 ;
wire \Add0~40_combout ;
wire \Add0~43 ;
wire \Add0~42_combout ;
wire \Add0~45 ;
wire \Add0~44_combout ;
wire \Add0~47 ;
wire \Add0~46_combout ;
wire \Add0~49 ;
wire \Add0~48_combout ;
wire \Add0~51 ;
wire \Add0~50_combout ;
wire \Add0~53 ;
wire \Add0~52_combout ;
wire \Add0~55 ;
wire \Add0~54_combout ;
wire \Add0~57 ;
wire \Add0~56_combout ;
wire \Add0~58_combout ;
wire \CU|Equal6~1_combout ;
wire \RF|Mux30~9_combout ;
wire \RF|Mux30~19_combout ;
wire \RF|Mux30~20_combout ;
wire \CU|Equal0~2_combout ;
wire \CU|always0~1_combout ;
wire \CU|cuif.RegWEN~0_combout ;
wire \CU|Equal7~0_combout ;
wire \CU|Equal3~0_combout ;
wire \CU|cuif.ALUOP[3]~8_combout ;
wire \CU|cuif.ALUOP[2]~11_combout ;
wire \CU|cuif.ALUOP[1]~16_combout ;
wire \CU|cuif.ALUOP[0]~19_combout ;
wire \RF|Mux0~20_combout ;
wire \portB~0_combout ;
wire \portB~1_combout ;
wire \portB~2_combout ;
wire \portB~3_combout ;
wire \RF|Mux1~20_combout ;
wire \portB~4_combout ;
wire \portB~5_combout ;
wire \RF|Mux2~20_combout ;
wire \portB~6_combout ;
wire \portB~7_combout ;
wire \RF|Mux3~20_combout ;
wire \portB~8_combout ;
wire \portB~9_combout ;
wire \RF|Mux4~20_combout ;
wire \portB~10_combout ;
wire \portB~11_combout ;
wire \RF|Mux5~20_combout ;
wire \portB~12_combout ;
wire \portB~13_combout ;
wire \RF|Mux6~20_combout ;
wire \portB~14_combout ;
wire \portB~15_combout ;
wire \RF|Mux7~9_combout ;
wire \RF|Mux7~19_combout ;
wire \RF|Mux7~20_combout ;
wire \portB~16_combout ;
wire \portB~17_combout ;
wire \RF|Mux8~20_combout ;
wire \portB~18_combout ;
wire \portB~19_combout ;
wire \RF|Mux9~20_combout ;
wire \portB~20_combout ;
wire \portB~21_combout ;
wire \RF|Mux10~20_combout ;
wire \portB~22_combout ;
wire \portB~23_combout ;
wire \RF|Mux11~20_combout ;
wire \portB~24_combout ;
wire \portB~25_combout ;
wire \RF|Mux12~20_combout ;
wire \portB~26_combout ;
wire \portB~27_combout ;
wire \RF|Mux13~20_combout ;
wire \portB~28_combout ;
wire \portB~29_combout ;
wire \RF|Mux14~20_combout ;
wire \portB~30_combout ;
wire \portB~31_combout ;
wire \RF|Mux15~20_combout ;
wire \portB~32_combout ;
wire \portB~33_combout ;
wire \RF|Mux16~20_combout ;
wire \portB~34_combout ;
wire \portB~35_combout ;
wire \RF|Mux17~20_combout ;
wire \portB~36_combout ;
wire \portB~37_combout ;
wire \RF|Mux18~20_combout ;
wire \portB~38_combout ;
wire \portB~39_combout ;
wire \RF|Mux19~20_combout ;
wire \portB~40_combout ;
wire \portB~41_combout ;
wire \RF|Mux20~20_combout ;
wire \portB~42_combout ;
wire \portB~43_combout ;
wire \RF|Mux21~20_combout ;
wire \portB~44_combout ;
wire \portB~45_combout ;
wire \RF|Mux22~20_combout ;
wire \portB~46_combout ;
wire \portB~47_combout ;
wire \RF|Mux23~20_combout ;
wire \portB~48_combout ;
wire \portB~49_combout ;
wire \RF|Mux24~9_combout ;
wire \RF|Mux24~19_combout ;
wire \RF|Mux24~20_combout ;
wire \portB~50_combout ;
wire \portB~51_combout ;
wire \RF|Mux25~9_combout ;
wire \RF|Mux25~19_combout ;
wire \RF|Mux25~20_combout ;
wire \portB~52_combout ;
wire \portB~53_combout ;
wire \RF|Mux26~20_combout ;
wire \portB~54_combout ;
wire \portB~55_combout ;
wire \RF|Mux27~9_combout ;
wire \RF|Mux27~19_combout ;
wire \RF|Mux27~20_combout ;
wire \portB~56_combout ;
wire \portB~57_combout ;
wire \RF|Mux28~20_combout ;
wire \portB~58_combout ;
wire \portB~59_combout ;
wire \RF|Mux29~9_combout ;
wire \RF|Mux29~19_combout ;
wire \RF|Mux29~20_combout ;
wire \portB~60_combout ;
wire \portB~61_combout ;
wire \portB~62_combout ;
wire \portB~63_combout ;
wire \RF|Mux31~9_combout ;
wire \RF|Mux31~19_combout ;
wire \RF|Mux31~20_combout ;
wire \portB~64_combout ;
wire \portB~65_combout ;
wire \ALU|Selector11~9_combout ;
wire \ALU|Selector29~8_combout ;
wire \ALU|Selector10~8_combout ;
wire \ALU|Selector5~8_combout ;
wire \ALU|Selector14~8_combout ;
wire \ALU|Selector26~8_combout ;
wire \ALU|Selector21~8_combout ;
wire \ALU|Selector8~10_combout ;
wire \ALU|Selector9~8_combout ;
wire \ALU|Equal0~11_combout ;
wire \CU|Equal2~2_combout ;
wire \CU|Equal3~1_combout ;
wire \CU|cuif.PCSrc[0]~1_combout ;
wire \CU|cuif.PCSrc[1]~2_combout ;
wire \CU|cuif.MemtoReg[0]~0_combout ;
wire \CU|cuif.MemtoReg[1]~1_combout ;
wire \wdat~0_combout ;
wire \wdat~1_combout ;
wire \CU|cuif.RegWEN~2_combout ;
wire \wsel~0_combout ;
wire \wsel~1_combout ;
wire \wsel~2_combout ;
wire \wsel~3_combout ;
wire \wsel~4_combout ;
wire \wdat~2_combout ;
wire \wdat~3_combout ;
wire \wdat~4_combout ;
wire \wdat~5_combout ;
wire \wdat~6_combout ;
wire \wdat~7_combout ;
wire \wdat~8_combout ;
wire \wdat~9_combout ;
wire \wdat~10_combout ;
wire \wdat~11_combout ;
wire \wdat~12_combout ;
wire \wdat~13_combout ;
wire \wdat~14_combout ;
wire \wdat~15_combout ;
wire \wdat~16_combout ;
wire \wdat~17_combout ;
wire \wdat~18_combout ;
wire \wdat~19_combout ;
wire \wdat~20_combout ;
wire \wdat~21_combout ;
wire \wdat~22_combout ;
wire \wdat~23_combout ;
wire \wdat~24_combout ;
wire \wdat~25_combout ;
wire \wdat~26_combout ;
wire \wdat~27_combout ;
wire \wdat~28_combout ;
wire \wdat~29_combout ;
wire \wdat~30_combout ;
wire \wdat~31_combout ;
wire \wdat~32_combout ;
wire \wdat~33_combout ;
wire \wdat~34_combout ;
wire \wdat~35_combout ;
wire \wdat~36_combout ;
wire \wdat~37_combout ;
wire \wdat~38_combout ;
wire \wdat~39_combout ;
wire \wdat~40_combout ;
wire \wdat~41_combout ;
wire \wdat~42_combout ;
wire \wdat~43_combout ;
wire \wdat~44_combout ;
wire \ALU|Selector20~9_combout ;
wire \wdat~45_combout ;
wire \wdat~46_combout ;
wire \wdat~47_combout ;
wire \wdat~48_combout ;
wire \wdat~49_combout ;
wire \wdat~50_combout ;
wire \wdat~51_combout ;
wire \wdat~52_combout ;
wire \wdat~53_combout ;
wire \wdat~54_combout ;
wire \wdat~55_combout ;
wire \wdat~56_combout ;
wire \wdat~57_combout ;
wire \wdat~58_combout ;
wire \wdat~59_combout ;
wire \wdat~60_combout ;
wire \wdat~61_combout ;
wire \wdat~62_combout ;
wire \wdat~63_combout ;
wire \CU|cuif.ALUOP[2]~20_combout ;
wire \ALU|Selector31~12_combout ;
wire \ALU|Selector23~11_combout ;


register_file RF(
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ccifiwait_0(ccifiwait_0),
	.dcifimemload_19(dcifimemload_19),
	.dcifimemload_18(dcifimemload_18),
	.instr_16(instr_16),
	.dcifimemload_16(dcifimemload_16),
	.instr_17(instr_17),
	.dcifimemload_17(dcifimemload_17),
	.Mux63(Mux63),
	.Mux631(Mux631),
	.dcifimemload_24(dcifimemload_24),
	.dcifimemload_23(dcifimemload_23),
	.dcifimemload_21(dcifimemload_21),
	.dcifimemload_22(dcifimemload_22),
	.Mux30(\RF|Mux30~9_combout ),
	.Mux301(\RF|Mux30~19_combout ),
	.dcifimemload_25(dcifimemload_25),
	.Mux302(\RF|Mux30~20_combout ),
	.Mux0(\RF|Mux0~20_combout ),
	.Mux32(Mux32),
	.Mux321(Mux321),
	.Mux1(\RF|Mux1~20_combout ),
	.Mux33(Mux33),
	.Mux331(Mux331),
	.Mux2(\RF|Mux2~20_combout ),
	.Mux34(Mux34),
	.Mux341(Mux341),
	.Mux3(\RF|Mux3~20_combout ),
	.Mux35(Mux35),
	.Mux351(Mux351),
	.Mux4(\RF|Mux4~20_combout ),
	.Mux36(Mux36),
	.Mux361(Mux361),
	.Mux5(\RF|Mux5~20_combout ),
	.Mux37(Mux37),
	.Mux371(Mux371),
	.Mux6(\RF|Mux6~20_combout ),
	.Mux38(Mux38),
	.Mux381(Mux381),
	.Mux7(\RF|Mux7~9_combout ),
	.Mux71(\RF|Mux7~19_combout ),
	.Mux72(\RF|Mux7~20_combout ),
	.Mux39(Mux39),
	.Mux391(Mux391),
	.Mux8(\RF|Mux8~20_combout ),
	.Mux40(Mux40),
	.Mux401(Mux401),
	.Mux9(\RF|Mux9~20_combout ),
	.Mux41(Mux41),
	.Mux411(Mux411),
	.Mux10(\RF|Mux10~20_combout ),
	.Mux42(Mux42),
	.Mux421(Mux421),
	.Mux11(\RF|Mux11~20_combout ),
	.Mux43(Mux43),
	.Mux431(Mux431),
	.Mux12(\RF|Mux12~20_combout ),
	.Mux44(Mux44),
	.Mux441(Mux441),
	.Mux13(\RF|Mux13~20_combout ),
	.Mux45(Mux45),
	.Mux451(Mux451),
	.Mux14(\RF|Mux14~20_combout ),
	.Mux46(Mux46),
	.Mux461(Mux461),
	.Mux15(\RF|Mux15~20_combout ),
	.Mux47(Mux47),
	.Mux471(Mux471),
	.Mux16(\RF|Mux16~20_combout ),
	.Mux48(Mux48),
	.Mux481(Mux481),
	.Mux17(\RF|Mux17~20_combout ),
	.Mux49(Mux49),
	.Mux491(Mux491),
	.Mux18(\RF|Mux18~20_combout ),
	.Mux50(Mux50),
	.Mux501(Mux501),
	.Mux19(\RF|Mux19~20_combout ),
	.Mux51(Mux51),
	.Mux511(Mux511),
	.Mux20(\RF|Mux20~20_combout ),
	.Mux52(Mux52),
	.Mux521(Mux521),
	.Mux21(\RF|Mux21~20_combout ),
	.Mux53(Mux53),
	.Mux531(Mux531),
	.Mux22(\RF|Mux22~20_combout ),
	.Mux54(Mux54),
	.Mux541(Mux541),
	.Mux23(\RF|Mux23~20_combout ),
	.Mux55(Mux55),
	.Mux551(Mux551),
	.Mux24(\RF|Mux24~9_combout ),
	.Mux241(\RF|Mux24~19_combout ),
	.Mux242(\RF|Mux24~20_combout ),
	.Mux56(Mux56),
	.Mux561(Mux561),
	.Mux25(\RF|Mux25~9_combout ),
	.Mux251(\RF|Mux25~19_combout ),
	.Mux252(\RF|Mux25~20_combout ),
	.Mux57(Mux57),
	.Mux571(Mux571),
	.Mux26(\RF|Mux26~20_combout ),
	.Mux58(Mux58),
	.Mux581(Mux581),
	.Mux27(\RF|Mux27~9_combout ),
	.Mux271(\RF|Mux27~19_combout ),
	.Mux272(\RF|Mux27~20_combout ),
	.Mux59(Mux59),
	.Mux591(Mux591),
	.Mux28(\RF|Mux28~20_combout ),
	.Mux60(Mux60),
	.Mux601(Mux601),
	.Mux29(\RF|Mux29~9_combout ),
	.Mux291(\RF|Mux29~19_combout ),
	.Mux292(\RF|Mux29~20_combout ),
	.Mux61(Mux61),
	.Mux611(Mux611),
	.Mux62(Mux62),
	.Mux621(Mux621),
	.Mux31(\RF|Mux31~9_combout ),
	.Mux311(\RF|Mux31~19_combout ),
	.Mux312(\RF|Mux31~20_combout ),
	.wdat(\wdat~1_combout ),
	.cuifRegWEN(\CU|cuif.RegWEN~2_combout ),
	.wsel(\wsel~0_combout ),
	.wsel1(\wsel~1_combout ),
	.wsel2(\wsel~2_combout ),
	.wsel3(\wsel~3_combout ),
	.wsel4(\wsel~4_combout ),
	.wdat1(\wdat~3_combout ),
	.wdat2(\wdat~5_combout ),
	.wdat3(\wdat~7_combout ),
	.wdat4(\wdat~9_combout ),
	.wdat5(\wdat~11_combout ),
	.wdat6(\wdat~13_combout ),
	.wdat7(\wdat~15_combout ),
	.wdat8(\wdat~17_combout ),
	.wdat9(\wdat~19_combout ),
	.wdat10(\wdat~21_combout ),
	.wdat11(\wdat~23_combout ),
	.wdat12(\wdat~25_combout ),
	.wdat13(\wdat~27_combout ),
	.wdat14(\wdat~29_combout ),
	.wdat15(\wdat~31_combout ),
	.wdat16(\wdat~33_combout ),
	.wdat17(\wdat~35_combout ),
	.wdat18(\wdat~37_combout ),
	.wdat19(\wdat~39_combout ),
	.wdat20(\wdat~41_combout ),
	.wdat21(\wdat~43_combout ),
	.wdat22(\wdat~45_combout ),
	.wdat23(\wdat~47_combout ),
	.wdat24(\wdat~49_combout ),
	.wdat25(\wdat~51_combout ),
	.wdat26(\wdat~53_combout ),
	.wdat27(\wdat~55_combout ),
	.wdat28(\wdat~57_combout ),
	.wdat29(\wdat~59_combout ),
	.wdat30(\wdat~61_combout ),
	.wdat31(\wdat~63_combout ),
	.CLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

alu ALU(
	.Mux30(\RF|Mux30~9_combout ),
	.Mux301(\RF|Mux30~19_combout ),
	.dcifimemload_25(dcifimemload_25),
	.Mux302(\RF|Mux30~20_combout ),
	.cuifALUOP_3(\CU|cuif.ALUOP[3]~8_combout ),
	.cuifALUOP_2(\CU|cuif.ALUOP[2]~11_combout ),
	.cuifALUOP_1(\CU|cuif.ALUOP[1]~16_combout ),
	.cuifALUOP_0(\CU|cuif.ALUOP[0]~19_combout ),
	.Mux0(\RF|Mux0~20_combout ),
	.portB(\portB~3_combout ),
	.Mux1(\RF|Mux1~20_combout ),
	.portB1(\portB~5_combout ),
	.Mux2(\RF|Mux2~20_combout ),
	.portB2(\portB~7_combout ),
	.Mux3(\RF|Mux3~20_combout ),
	.portB3(\portB~9_combout ),
	.Mux4(\RF|Mux4~20_combout ),
	.portB4(\portB~11_combout ),
	.Mux5(\RF|Mux5~20_combout ),
	.portB5(\portB~13_combout ),
	.Mux6(\RF|Mux6~20_combout ),
	.portB6(\portB~15_combout ),
	.Mux7(\RF|Mux7~9_combout ),
	.Mux71(\RF|Mux7~19_combout ),
	.Mux72(\RF|Mux7~20_combout ),
	.portB7(\portB~17_combout ),
	.Mux8(\RF|Mux8~20_combout ),
	.portB8(\portB~19_combout ),
	.Mux9(\RF|Mux9~20_combout ),
	.portB9(\portB~21_combout ),
	.Mux10(\RF|Mux10~20_combout ),
	.portB10(\portB~23_combout ),
	.Mux11(\RF|Mux11~20_combout ),
	.portB11(\portB~25_combout ),
	.Mux12(\RF|Mux12~20_combout ),
	.portB12(\portB~27_combout ),
	.Mux13(\RF|Mux13~20_combout ),
	.portB13(\portB~29_combout ),
	.Mux14(\RF|Mux14~20_combout ),
	.portB14(\portB~31_combout ),
	.Mux15(\RF|Mux15~20_combout ),
	.portB15(\portB~33_combout ),
	.Mux16(\RF|Mux16~20_combout ),
	.portB16(\portB~35_combout ),
	.Mux17(\RF|Mux17~20_combout ),
	.portB17(\portB~37_combout ),
	.Mux18(\RF|Mux18~20_combout ),
	.portB18(\portB~39_combout ),
	.Mux19(\RF|Mux19~20_combout ),
	.portB19(\portB~41_combout ),
	.Mux20(\RF|Mux20~20_combout ),
	.portB20(\portB~43_combout ),
	.Mux21(\RF|Mux21~20_combout ),
	.portB21(\portB~45_combout ),
	.Mux22(\RF|Mux22~20_combout ),
	.portB22(\portB~47_combout ),
	.Mux23(\RF|Mux23~20_combout ),
	.portB23(\portB~49_combout ),
	.Mux24(\RF|Mux24~9_combout ),
	.Mux241(\RF|Mux24~19_combout ),
	.Mux242(\RF|Mux24~20_combout ),
	.portB24(\portB~51_combout ),
	.Mux25(\RF|Mux25~9_combout ),
	.Mux251(\RF|Mux25~19_combout ),
	.Mux252(\RF|Mux25~20_combout ),
	.portB25(\portB~53_combout ),
	.Mux26(\RF|Mux26~20_combout ),
	.portB26(\portB~55_combout ),
	.Mux27(\RF|Mux27~9_combout ),
	.Mux271(\RF|Mux27~19_combout ),
	.Mux272(\RF|Mux27~20_combout ),
	.portB27(\portB~57_combout ),
	.Mux28(\RF|Mux28~20_combout ),
	.portB28(\portB~59_combout ),
	.Mux29(\RF|Mux29~9_combout ),
	.Mux291(\RF|Mux29~19_combout ),
	.Mux292(\RF|Mux29~20_combout ),
	.portB29(\portB~61_combout ),
	.portB30(\portB~63_combout ),
	.Mux31(\RF|Mux31~9_combout ),
	.Mux311(\RF|Mux31~19_combout ),
	.Mux312(\RF|Mux31~20_combout ),
	.portB31(\portB~65_combout ),
	.Selector31(Selector31),
	.ShiftRight0(ShiftRight0),
	.Selector24(Selector24),
	.Selector8(Selector8),
	.Selector0(Selector0),
	.Selector3(Selector3),
	.Selector4(Selector4),
	.Selector7(Selector7),
	.Selector11(Selector11),
	.ShiftRight01(ShiftRight01),
	.Selector111(\ALU|Selector11~9_combout ),
	.Selector15(Selector15),
	.Selector22(Selector22),
	.Selector28(Selector28),
	.Selector29(Selector29),
	.ShiftRight02(ShiftRight02),
	.ShiftRight03(ShiftRight03),
	.Selector291(\ALU|Selector29~8_combout ),
	.ShiftLeft0(ShiftLeft0),
	.Selector10(Selector10),
	.Selector101(Selector101),
	.Selector102(Selector102),
	.Selector103(\ALU|Selector10~8_combout ),
	.Selector2(Selector2),
	.Selector1(Selector1),
	.Selector41(Selector41),
	.Selector5(Selector5),
	.Selector51(\ALU|Selector5~8_combout ),
	.Selector12(Selector12),
	.Selector241(Selector241),
	.Selector242(Selector242),
	.Selector13(Selector13),
	.Selector25(Selector25),
	.Selector14(Selector14),
	.Selector141(Selector141),
	.Selector142(Selector142),
	.Selector143(\ALU|Selector14~8_combout ),
	.Selector27(Selector27),
	.Selector16(Selector16),
	.Selector18(Selector18),
	.Selector17(Selector17),
	.Selector6(Selector6),
	.Selector26(Selector26),
	.Selector261(\ALU|Selector26~8_combout ),
	.Selector19(Selector19),
	.Selector20(Selector20),
	.Selector201(Selector201),
	.Selector202(Selector202),
	.Selector21(Selector21),
	.Selector211(Selector211),
	.Selector212(Selector212),
	.Selector213(\ALU|Selector21~8_combout ),
	.Selector81(Selector81),
	.Selector82(Selector82),
	.Selector83(Selector83),
	.Selector84(\ALU|Selector8~10_combout ),
	.Selector9(Selector9),
	.Selector91(Selector91),
	.Selector92(Selector92),
	.Selector93(\ALU|Selector9~8_combout ),
	.Selector221(Selector221),
	.Selector30(Selector30),
	.Selector23(Selector23),
	.Selector231(Selector231),
	.Selector232(Selector232),
	.Equal0(\ALU|Equal0~11_combout ),
	.Selector203(\ALU|Selector20~9_combout ),
	.Selector311(\ALU|Selector31~12_combout ),
	.Selector233(\ALU|Selector23~11_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

control_unit CU(
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.instr_30(instr_30),
	.ccifiwait_0(ccifiwait_0),
	.dcifimemload_30(dcifimemload_30),
	.instr_31(instr_31),
	.dcifimemload_31(dcifimemload_31),
	.instr_27(instr_27),
	.dcifimemload_27(dcifimemload_27),
	.instr_26(instr_26),
	.dcifimemload_26(dcifimemload_26),
	.instr_29(instr_29),
	.dcifimemload_29(dcifimemload_29),
	.instr_28(instr_28),
	.dcifimemload_28(dcifimemload_28),
	.Equal6(\CU|Equal6~1_combout ),
	.Equal0(\CU|Equal0~2_combout ),
	.dcifimemload_3(dcifimemload_3),
	.dcifimemload_4(dcifimemload_4),
	.dcifimemload_2(dcifimemload_2),
	.dcifimemload_5(dcifimemload_5),
	.dcifimemload_0(dcifimemload_0),
	.dcifimemload_1(dcifimemload_1),
	.always0(\CU|always0~1_combout ),
	.cuifRegWEN(\CU|cuif.RegWEN~0_combout ),
	.Equal7(\CU|Equal7~0_combout ),
	.Equal3(\CU|Equal3~0_combout ),
	.cuifALUOP_3(\CU|cuif.ALUOP[3]~8_combout ),
	.cuifALUOP_2(\CU|cuif.ALUOP[2]~11_combout ),
	.cuifALUOP_1(\CU|cuif.ALUOP[1]~16_combout ),
	.cuifALUOP_0(\CU|cuif.ALUOP[0]~19_combout ),
	.Equal01(\ALU|Equal0~11_combout ),
	.Equal2(\CU|Equal2~2_combout ),
	.Equal31(\CU|Equal3~1_combout ),
	.cuifPCSrc_0(\CU|cuif.PCSrc[0]~1_combout ),
	.dcifdhit(dcifdhit),
	.cuifPCSrc_1(\CU|cuif.PCSrc[1]~2_combout ),
	.cuifMemtoReg_0(\CU|cuif.MemtoReg[0]~0_combout ),
	.cuifMemtoReg_1(\CU|cuif.MemtoReg[1]~1_combout ),
	.cuifRegWEN1(\CU|cuif.RegWEN~2_combout ),
	.cuifALUOP_21(\CU|cuif.ALUOP[2]~20_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

request_unit RU(
	.reg_WEN1(reg_WEN),
	.reg_REN1(reg_REN),
	.always1(always1),
	.dcifimemload_31(dcifimemload_31),
	.dcifimemload_29(dcifimemload_29),
	.Equal3(\CU|Equal3~0_combout ),
	.dcifdhit(dcifdhit),
	.CLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

program_counter_unit PCU(
	.PC_29(PC_29),
	.PC_28(PC_28),
	.PC_31(PC_31),
	.PC_30(PC_30),
	.PC_1(PC_1),
	.PC_0(PC_0),
	.PC_3(PC_3),
	.PC_2(PC_2),
	.PC_5(PC_5),
	.PC_4(PC_4),
	.PC_7(PC_7),
	.PC_6(PC_6),
	.PC_9(PC_9),
	.PC_8(PC_8),
	.PC_11(PC_11),
	.PC_10(PC_10),
	.PC_13(PC_13),
	.PC_12(PC_12),
	.PC_15(PC_15),
	.PC_14(PC_14),
	.PC_17(PC_17),
	.PC_16(PC_16),
	.PC_19(PC_19),
	.PC_18(PC_18),
	.PC_21(PC_21),
	.PC_20(PC_20),
	.PC_23(PC_23),
	.PC_22(PC_22),
	.PC_25(PC_25),
	.PC_24(PC_24),
	.PC_27(PC_27),
	.PC_26(PC_26),
	.\pcuif.ihit (ccifiwait_0),
	.dcifimemload_19(dcifimemload_19),
	.dcifimemload_18(dcifimemload_18),
	.dcifimemload_16(dcifimemload_16),
	.dcifimemload_17(dcifimemload_17),
	.dcifimemload_20(dcifimemload_20),
	.dcifimemload_24(dcifimemload_24),
	.dcifimemload_23(dcifimemload_23),
	.dcifimemload_21(dcifimemload_21),
	.dcifimemload_22(dcifimemload_22),
	.Mux30(\RF|Mux30~9_combout ),
	.Mux301(\RF|Mux30~19_combout ),
	.dcifimemload_25(dcifimemload_25),
	.dcifimemload_3(dcifimemload_3),
	.dcifimemload_4(dcifimemload_4),
	.dcifimemload_2(dcifimemload_2),
	.dcifimemload_5(dcifimemload_5),
	.dcifimemload_0(dcifimemload_0),
	.dcifimemload_1(dcifimemload_1),
	.always0(\CU|always0~1_combout ),
	.Mux0(\RF|Mux0~20_combout ),
	.dcifimemload_15(dcifimemload_15),
	.Mux1(\RF|Mux1~20_combout ),
	.Mux2(\RF|Mux2~20_combout ),
	.Mux3(\RF|Mux3~20_combout ),
	.Mux4(\RF|Mux4~20_combout ),
	.Mux5(\RF|Mux5~20_combout ),
	.Mux6(\RF|Mux6~20_combout ),
	.Mux7(\RF|Mux7~20_combout ),
	.Mux8(\RF|Mux8~20_combout ),
	.Mux9(\RF|Mux9~20_combout ),
	.Mux10(\RF|Mux10~20_combout ),
	.Mux11(\RF|Mux11~20_combout ),
	.Mux12(\RF|Mux12~20_combout ),
	.Mux13(\RF|Mux13~20_combout ),
	.Mux14(\RF|Mux14~20_combout ),
	.Mux15(\RF|Mux15~20_combout ),
	.Mux16(\RF|Mux16~20_combout ),
	.Mux17(\RF|Mux17~20_combout ),
	.dcifimemload_14(dcifimemload_14),
	.Mux18(\RF|Mux18~20_combout ),
	.dcifimemload_13(dcifimemload_13),
	.Mux19(\RF|Mux19~20_combout ),
	.dcifimemload_12(dcifimemload_12),
	.Mux20(\RF|Mux20~20_combout ),
	.dcifimemload_11(dcifimemload_11),
	.Mux21(\RF|Mux21~20_combout ),
	.dcifimemload_10(dcifimemload_10),
	.Mux22(\RF|Mux22~20_combout ),
	.dcifimemload_9(dcifimemload_9),
	.Mux23(\RF|Mux23~20_combout ),
	.dcifimemload_8(dcifimemload_8),
	.Mux24(\RF|Mux24~20_combout ),
	.dcifimemload_7(dcifimemload_7),
	.Mux25(\RF|Mux25~20_combout ),
	.dcifimemload_6(dcifimemload_6),
	.Mux26(\RF|Mux26~20_combout ),
	.Mux27(\RF|Mux27~20_combout ),
	.Mux28(\RF|Mux28~20_combout ),
	.Mux29(\RF|Mux29~20_combout ),
	.Mux31(\RF|Mux31~9_combout ),
	.Mux311(\RF|Mux31~19_combout ),
	.Equal2(\CU|Equal2~2_combout ),
	.Equal3(\CU|Equal3~1_combout ),
	.cuifPCSrc_0(\CU|cuif.PCSrc[0]~1_combout ),
	.cuifPCSrc_1(\CU|cuif.PCSrc[1]~2_combout ),
	.CLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X58_Y29_N2
cycloneive_lcell_comb \Add0~0 (
// Equation(s):
// \Add0~0_combout  = PC_2 $ (VCC)
// \Add0~1  = CARRY(PC_2)

	.dataa(gnd),
	.datab(PC_2),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
// synopsys translate_off
defparam \Add0~0 .lut_mask = 16'h33CC;
defparam \Add0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N4
cycloneive_lcell_comb \Add0~2 (
// Equation(s):
// \Add0~2_combout  = (PC_3 & (!\Add0~1 )) # (!PC_3 & ((\Add0~1 ) # (GND)))
// \Add0~3  = CARRY((!\Add0~1 ) # (!PC_3))

	.dataa(gnd),
	.datab(PC_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
// synopsys translate_off
defparam \Add0~2 .lut_mask = 16'h3C3F;
defparam \Add0~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N6
cycloneive_lcell_comb \Add0~4 (
// Equation(s):
// \Add0~4_combout  = (PC_4 & (\Add0~3  $ (GND))) # (!PC_4 & (!\Add0~3  & VCC))
// \Add0~5  = CARRY((PC_4 & !\Add0~3 ))

	.dataa(gnd),
	.datab(PC_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
// synopsys translate_off
defparam \Add0~4 .lut_mask = 16'hC30C;
defparam \Add0~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N8
cycloneive_lcell_comb \Add0~6 (
// Equation(s):
// \Add0~6_combout  = (PC_5 & (!\Add0~5 )) # (!PC_5 & ((\Add0~5 ) # (GND)))
// \Add0~7  = CARRY((!\Add0~5 ) # (!PC_5))

	.dataa(gnd),
	.datab(PC_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
// synopsys translate_off
defparam \Add0~6 .lut_mask = 16'h3C3F;
defparam \Add0~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N10
cycloneive_lcell_comb \Add0~8 (
// Equation(s):
// \Add0~8_combout  = (PC_6 & (\Add0~7  $ (GND))) # (!PC_6 & (!\Add0~7  & VCC))
// \Add0~9  = CARRY((PC_6 & !\Add0~7 ))

	.dataa(gnd),
	.datab(PC_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
// synopsys translate_off
defparam \Add0~8 .lut_mask = 16'hC30C;
defparam \Add0~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N12
cycloneive_lcell_comb \Add0~10 (
// Equation(s):
// \Add0~10_combout  = (PC_7 & (!\Add0~9 )) # (!PC_7 & ((\Add0~9 ) # (GND)))
// \Add0~11  = CARRY((!\Add0~9 ) # (!PC_7))

	.dataa(gnd),
	.datab(PC_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
// synopsys translate_off
defparam \Add0~10 .lut_mask = 16'h3C3F;
defparam \Add0~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N14
cycloneive_lcell_comb \Add0~12 (
// Equation(s):
// \Add0~12_combout  = (PC_8 & (\Add0~11  $ (GND))) # (!PC_8 & (!\Add0~11  & VCC))
// \Add0~13  = CARRY((PC_8 & !\Add0~11 ))

	.dataa(gnd),
	.datab(PC_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
// synopsys translate_off
defparam \Add0~12 .lut_mask = 16'hC30C;
defparam \Add0~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N16
cycloneive_lcell_comb \Add0~14 (
// Equation(s):
// \Add0~14_combout  = (PC_9 & (!\Add0~13 )) # (!PC_9 & ((\Add0~13 ) # (GND)))
// \Add0~15  = CARRY((!\Add0~13 ) # (!PC_9))

	.dataa(PC_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
// synopsys translate_off
defparam \Add0~14 .lut_mask = 16'h5A5F;
defparam \Add0~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N18
cycloneive_lcell_comb \Add0~16 (
// Equation(s):
// \Add0~16_combout  = (PC_10 & (\Add0~15  $ (GND))) # (!PC_10 & (!\Add0~15  & VCC))
// \Add0~17  = CARRY((PC_10 & !\Add0~15 ))

	.dataa(gnd),
	.datab(PC_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
// synopsys translate_off
defparam \Add0~16 .lut_mask = 16'hC30C;
defparam \Add0~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N20
cycloneive_lcell_comb \Add0~18 (
// Equation(s):
// \Add0~18_combout  = (PC_11 & (!\Add0~17 )) # (!PC_11 & ((\Add0~17 ) # (GND)))
// \Add0~19  = CARRY((!\Add0~17 ) # (!PC_11))

	.dataa(gnd),
	.datab(PC_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
// synopsys translate_off
defparam \Add0~18 .lut_mask = 16'h3C3F;
defparam \Add0~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N22
cycloneive_lcell_comb \Add0~20 (
// Equation(s):
// \Add0~20_combout  = (PC_12 & (\Add0~19  $ (GND))) # (!PC_12 & (!\Add0~19  & VCC))
// \Add0~21  = CARRY((PC_12 & !\Add0~19 ))

	.dataa(PC_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
// synopsys translate_off
defparam \Add0~20 .lut_mask = 16'hA50A;
defparam \Add0~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N24
cycloneive_lcell_comb \Add0~22 (
// Equation(s):
// \Add0~22_combout  = (PC_13 & (!\Add0~21 )) # (!PC_13 & ((\Add0~21 ) # (GND)))
// \Add0~23  = CARRY((!\Add0~21 ) # (!PC_13))

	.dataa(PC_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
// synopsys translate_off
defparam \Add0~22 .lut_mask = 16'h5A5F;
defparam \Add0~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N26
cycloneive_lcell_comb \Add0~24 (
// Equation(s):
// \Add0~24_combout  = (PC_14 & (\Add0~23  $ (GND))) # (!PC_14 & (!\Add0~23  & VCC))
// \Add0~25  = CARRY((PC_14 & !\Add0~23 ))

	.dataa(PC_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
// synopsys translate_off
defparam \Add0~24 .lut_mask = 16'hA50A;
defparam \Add0~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N28
cycloneive_lcell_comb \Add0~26 (
// Equation(s):
// \Add0~26_combout  = (PC_15 & (!\Add0~25 )) # (!PC_15 & ((\Add0~25 ) # (GND)))
// \Add0~27  = CARRY((!\Add0~25 ) # (!PC_15))

	.dataa(gnd),
	.datab(PC_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout(\Add0~27 ));
// synopsys translate_off
defparam \Add0~26 .lut_mask = 16'h3C3F;
defparam \Add0~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N30
cycloneive_lcell_comb \Add0~28 (
// Equation(s):
// \Add0~28_combout  = (PC_16 & (\Add0~27  $ (GND))) # (!PC_16 & (!\Add0~27  & VCC))
// \Add0~29  = CARRY((PC_16 & !\Add0~27 ))

	.dataa(PC_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~27 ),
	.combout(\Add0~28_combout ),
	.cout(\Add0~29 ));
// synopsys translate_off
defparam \Add0~28 .lut_mask = 16'hA50A;
defparam \Add0~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N0
cycloneive_lcell_comb \Add0~30 (
// Equation(s):
// \Add0~30_combout  = (PC_17 & (!\Add0~29 )) # (!PC_17 & ((\Add0~29 ) # (GND)))
// \Add0~31  = CARRY((!\Add0~29 ) # (!PC_17))

	.dataa(gnd),
	.datab(PC_17),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~29 ),
	.combout(\Add0~30_combout ),
	.cout(\Add0~31 ));
// synopsys translate_off
defparam \Add0~30 .lut_mask = 16'h3C3F;
defparam \Add0~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N2
cycloneive_lcell_comb \Add0~32 (
// Equation(s):
// \Add0~32_combout  = (PC_18 & (\Add0~31  $ (GND))) # (!PC_18 & (!\Add0~31  & VCC))
// \Add0~33  = CARRY((PC_18 & !\Add0~31 ))

	.dataa(PC_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~31 ),
	.combout(\Add0~32_combout ),
	.cout(\Add0~33 ));
// synopsys translate_off
defparam \Add0~32 .lut_mask = 16'hA50A;
defparam \Add0~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N4
cycloneive_lcell_comb \Add0~34 (
// Equation(s):
// \Add0~34_combout  = (PC_19 & (!\Add0~33 )) # (!PC_19 & ((\Add0~33 ) # (GND)))
// \Add0~35  = CARRY((!\Add0~33 ) # (!PC_19))

	.dataa(PC_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~33 ),
	.combout(\Add0~34_combout ),
	.cout(\Add0~35 ));
// synopsys translate_off
defparam \Add0~34 .lut_mask = 16'h5A5F;
defparam \Add0~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N6
cycloneive_lcell_comb \Add0~36 (
// Equation(s):
// \Add0~36_combout  = (PC_20 & (\Add0~35  $ (GND))) # (!PC_20 & (!\Add0~35  & VCC))
// \Add0~37  = CARRY((PC_20 & !\Add0~35 ))

	.dataa(PC_20),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~35 ),
	.combout(\Add0~36_combout ),
	.cout(\Add0~37 ));
// synopsys translate_off
defparam \Add0~36 .lut_mask = 16'hA50A;
defparam \Add0~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N8
cycloneive_lcell_comb \Add0~38 (
// Equation(s):
// \Add0~38_combout  = (PC_21 & (!\Add0~37 )) # (!PC_21 & ((\Add0~37 ) # (GND)))
// \Add0~39  = CARRY((!\Add0~37 ) # (!PC_21))

	.dataa(gnd),
	.datab(PC_21),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~37 ),
	.combout(\Add0~38_combout ),
	.cout(\Add0~39 ));
// synopsys translate_off
defparam \Add0~38 .lut_mask = 16'h3C3F;
defparam \Add0~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N10
cycloneive_lcell_comb \Add0~40 (
// Equation(s):
// \Add0~40_combout  = (PC_22 & (\Add0~39  $ (GND))) # (!PC_22 & (!\Add0~39  & VCC))
// \Add0~41  = CARRY((PC_22 & !\Add0~39 ))

	.dataa(PC_22),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~39 ),
	.combout(\Add0~40_combout ),
	.cout(\Add0~41 ));
// synopsys translate_off
defparam \Add0~40 .lut_mask = 16'hA50A;
defparam \Add0~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N12
cycloneive_lcell_comb \Add0~42 (
// Equation(s):
// \Add0~42_combout  = (PC_23 & (!\Add0~41 )) # (!PC_23 & ((\Add0~41 ) # (GND)))
// \Add0~43  = CARRY((!\Add0~41 ) # (!PC_23))

	.dataa(PC_23),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~41 ),
	.combout(\Add0~42_combout ),
	.cout(\Add0~43 ));
// synopsys translate_off
defparam \Add0~42 .lut_mask = 16'h5A5F;
defparam \Add0~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N14
cycloneive_lcell_comb \Add0~44 (
// Equation(s):
// \Add0~44_combout  = (PC_24 & (\Add0~43  $ (GND))) # (!PC_24 & (!\Add0~43  & VCC))
// \Add0~45  = CARRY((PC_24 & !\Add0~43 ))

	.dataa(PC_24),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~43 ),
	.combout(\Add0~44_combout ),
	.cout(\Add0~45 ));
// synopsys translate_off
defparam \Add0~44 .lut_mask = 16'hA50A;
defparam \Add0~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N16
cycloneive_lcell_comb \Add0~46 (
// Equation(s):
// \Add0~46_combout  = (PC_25 & (!\Add0~45 )) # (!PC_25 & ((\Add0~45 ) # (GND)))
// \Add0~47  = CARRY((!\Add0~45 ) # (!PC_25))

	.dataa(PC_25),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~45 ),
	.combout(\Add0~46_combout ),
	.cout(\Add0~47 ));
// synopsys translate_off
defparam \Add0~46 .lut_mask = 16'h5A5F;
defparam \Add0~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N18
cycloneive_lcell_comb \Add0~48 (
// Equation(s):
// \Add0~48_combout  = (PC_26 & (\Add0~47  $ (GND))) # (!PC_26 & (!\Add0~47  & VCC))
// \Add0~49  = CARRY((PC_26 & !\Add0~47 ))

	.dataa(gnd),
	.datab(PC_26),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~47 ),
	.combout(\Add0~48_combout ),
	.cout(\Add0~49 ));
// synopsys translate_off
defparam \Add0~48 .lut_mask = 16'hC30C;
defparam \Add0~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N20
cycloneive_lcell_comb \Add0~50 (
// Equation(s):
// \Add0~50_combout  = (PC_27 & (!\Add0~49 )) # (!PC_27 & ((\Add0~49 ) # (GND)))
// \Add0~51  = CARRY((!\Add0~49 ) # (!PC_27))

	.dataa(gnd),
	.datab(PC_27),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~49 ),
	.combout(\Add0~50_combout ),
	.cout(\Add0~51 ));
// synopsys translate_off
defparam \Add0~50 .lut_mask = 16'h3C3F;
defparam \Add0~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N22
cycloneive_lcell_comb \Add0~52 (
// Equation(s):
// \Add0~52_combout  = (PC_28 & (\Add0~51  $ (GND))) # (!PC_28 & (!\Add0~51  & VCC))
// \Add0~53  = CARRY((PC_28 & !\Add0~51 ))

	.dataa(PC_28),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~51 ),
	.combout(\Add0~52_combout ),
	.cout(\Add0~53 ));
// synopsys translate_off
defparam \Add0~52 .lut_mask = 16'hA50A;
defparam \Add0~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N24
cycloneive_lcell_comb \Add0~54 (
// Equation(s):
// \Add0~54_combout  = (PC_29 & (!\Add0~53 )) # (!PC_29 & ((\Add0~53 ) # (GND)))
// \Add0~55  = CARRY((!\Add0~53 ) # (!PC_29))

	.dataa(gnd),
	.datab(PC_29),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~53 ),
	.combout(\Add0~54_combout ),
	.cout(\Add0~55 ));
// synopsys translate_off
defparam \Add0~54 .lut_mask = 16'h3C3F;
defparam \Add0~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N26
cycloneive_lcell_comb \Add0~56 (
// Equation(s):
// \Add0~56_combout  = (PC_30 & (\Add0~55  $ (GND))) # (!PC_30 & (!\Add0~55  & VCC))
// \Add0~57  = CARRY((PC_30 & !\Add0~55 ))

	.dataa(gnd),
	.datab(PC_30),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~55 ),
	.combout(\Add0~56_combout ),
	.cout(\Add0~57 ));
// synopsys translate_off
defparam \Add0~56 .lut_mask = 16'hC30C;
defparam \Add0~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N28
cycloneive_lcell_comb \Add0~58 (
// Equation(s):
// \Add0~58_combout  = \Add0~57  $ (PC_31)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(PC_31),
	.cin(\Add0~57 ),
	.combout(\Add0~58_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~58 .lut_mask = 16'h0FF0;
defparam \Add0~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N6
cycloneive_lcell_comb \portB~0 (
// Equation(s):
// \portB~0_combout  = (dcifimemload_15 & (cuifRegWEN & !Equal0))

	.dataa(dcifimemload_15),
	.datab(gnd),
	.datac(\CU|cuif.RegWEN~0_combout ),
	.datad(\CU|Equal0~2_combout ),
	.cin(gnd),
	.combout(\portB~0_combout ),
	.cout());
// synopsys translate_off
defparam \portB~0 .lut_mask = 16'h00A0;
defparam \portB~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N28
cycloneive_lcell_comb \portB~1 (
// Equation(s):
// \portB~1_combout  = (\portB~0_combout  & (((dcifimemload_27 & dcifimemload_26)) # (!Equal7)))

	.dataa(\CU|Equal7~0_combout ),
	.datab(dcifimemload_27),
	.datac(dcifimemload_26),
	.datad(\portB~0_combout ),
	.cin(gnd),
	.combout(\portB~1_combout ),
	.cout());
// synopsys translate_off
defparam \portB~1 .lut_mask = 16'hD500;
defparam \portB~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N16
cycloneive_lcell_comb \portB~2 (
// Equation(s):
// \portB~2_combout  = (\portB~1_combout ) # ((Mux32 & (!cuifALUOP_21 & !dcifimemload_20)))

	.dataa(Mux32),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(dcifimemload_20),
	.datad(\portB~1_combout ),
	.cin(gnd),
	.combout(\portB~2_combout ),
	.cout());
// synopsys translate_off
defparam \portB~2 .lut_mask = 16'hFF02;
defparam \portB~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N22
cycloneive_lcell_comb \portB~3 (
// Equation(s):
// \portB~3_combout  = (\portB~2_combout ) # ((dcifimemload_20 & (Mux321 & !cuifALUOP_21)))

	.dataa(dcifimemload_20),
	.datab(Mux321),
	.datac(\CU|cuif.ALUOP[2]~20_combout ),
	.datad(\portB~2_combout ),
	.cin(gnd),
	.combout(\portB~3_combout ),
	.cout());
// synopsys translate_off
defparam \portB~3 .lut_mask = 16'hFF08;
defparam \portB~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N6
cycloneive_lcell_comb \portB~4 (
// Equation(s):
// \portB~4_combout  = (\portB~1_combout ) # ((!cuifALUOP_21 & (!dcifimemload_20 & Mux33)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(Mux33),
	.datad(\portB~1_combout ),
	.cin(gnd),
	.combout(\portB~4_combout ),
	.cout());
// synopsys translate_off
defparam \portB~4 .lut_mask = 16'hFF10;
defparam \portB~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N28
cycloneive_lcell_comb \portB~5 (
// Equation(s):
// \portB~5_combout  = (\portB~4_combout ) # ((Mux331 & (!cuifALUOP_21 & dcifimemload_20)))

	.dataa(Mux331),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(dcifimemload_20),
	.datad(\portB~4_combout ),
	.cin(gnd),
	.combout(\portB~5_combout ),
	.cout());
// synopsys translate_off
defparam \portB~5 .lut_mask = 16'hFF20;
defparam \portB~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N18
cycloneive_lcell_comb \portB~6 (
// Equation(s):
// \portB~6_combout  = (\portB~1_combout ) # ((!dcifimemload_20 & (!cuifALUOP_21 & Mux34)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(\portB~1_combout ),
	.datad(Mux34),
	.cin(gnd),
	.combout(\portB~6_combout ),
	.cout());
// synopsys translate_off
defparam \portB~6 .lut_mask = 16'hF1F0;
defparam \portB~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N26
cycloneive_lcell_comb \portB~7 (
// Equation(s):
// \portB~7_combout  = (\portB~6_combout ) # ((dcifimemload_20 & (!cuifALUOP_21 & Mux341)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux341),
	.datad(\portB~6_combout ),
	.cin(gnd),
	.combout(\portB~7_combout ),
	.cout());
// synopsys translate_off
defparam \portB~7 .lut_mask = 16'hFF20;
defparam \portB~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N24
cycloneive_lcell_comb \portB~8 (
// Equation(s):
// \portB~8_combout  = (\portB~1_combout ) # ((Mux35 & (!cuifALUOP_21 & !dcifimemload_20)))

	.dataa(Mux35),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(dcifimemload_20),
	.datad(\portB~1_combout ),
	.cin(gnd),
	.combout(\portB~8_combout ),
	.cout());
// synopsys translate_off
defparam \portB~8 .lut_mask = 16'hFF02;
defparam \portB~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N30
cycloneive_lcell_comb \portB~9 (
// Equation(s):
// \portB~9_combout  = (\portB~8_combout ) # ((dcifimemload_20 & (!cuifALUOP_21 & Mux351)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux351),
	.datad(\portB~8_combout ),
	.cin(gnd),
	.combout(\portB~9_combout ),
	.cout());
// synopsys translate_off
defparam \portB~9 .lut_mask = 16'hFF20;
defparam \portB~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N28
cycloneive_lcell_comb \portB~10 (
// Equation(s):
// \portB~10_combout  = (\portB~1_combout ) # ((!dcifimemload_20 & (!cuifALUOP_21 & Mux36)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux36),
	.datad(\portB~1_combout ),
	.cin(gnd),
	.combout(\portB~10_combout ),
	.cout());
// synopsys translate_off
defparam \portB~10 .lut_mask = 16'hFF10;
defparam \portB~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N18
cycloneive_lcell_comb \portB~11 (
// Equation(s):
// \portB~11_combout  = (\portB~10_combout ) # ((dcifimemload_20 & (!cuifALUOP_21 & Mux361)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux361),
	.datad(\portB~10_combout ),
	.cin(gnd),
	.combout(\portB~11_combout ),
	.cout());
// synopsys translate_off
defparam \portB~11 .lut_mask = 16'hFF20;
defparam \portB~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N12
cycloneive_lcell_comb \portB~12 (
// Equation(s):
// \portB~12_combout  = (\portB~1_combout ) # ((!cuifALUOP_21 & (!dcifimemload_20 & Mux37)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(Mux37),
	.datad(\portB~1_combout ),
	.cin(gnd),
	.combout(\portB~12_combout ),
	.cout());
// synopsys translate_off
defparam \portB~12 .lut_mask = 16'hFF10;
defparam \portB~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N10
cycloneive_lcell_comb \portB~13 (
// Equation(s):
// \portB~13_combout  = (\portB~12_combout ) # ((!cuifALUOP_21 & (dcifimemload_20 & Mux371)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(Mux371),
	.datad(\portB~12_combout ),
	.cin(gnd),
	.combout(\portB~13_combout ),
	.cout());
// synopsys translate_off
defparam \portB~13 .lut_mask = 16'hFF40;
defparam \portB~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N2
cycloneive_lcell_comb \portB~14 (
// Equation(s):
// \portB~14_combout  = (\portB~1_combout ) # ((!dcifimemload_20 & (!cuifALUOP_21 & Mux38)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(\portB~1_combout ),
	.datad(Mux38),
	.cin(gnd),
	.combout(\portB~14_combout ),
	.cout());
// synopsys translate_off
defparam \portB~14 .lut_mask = 16'hF1F0;
defparam \portB~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N4
cycloneive_lcell_comb \portB~15 (
// Equation(s):
// \portB~15_combout  = (\portB~14_combout ) # ((dcifimemload_20 & (!cuifALUOP_21 & Mux381)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux381),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~15_combout ),
	.cout());
// synopsys translate_off
defparam \portB~15 .lut_mask = 16'hFF20;
defparam \portB~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N26
cycloneive_lcell_comb \portB~16 (
// Equation(s):
// \portB~16_combout  = (\portB~1_combout ) # ((!dcifimemload_20 & (!cuifALUOP_21 & Mux39)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux39),
	.datad(\portB~1_combout ),
	.cin(gnd),
	.combout(\portB~16_combout ),
	.cout());
// synopsys translate_off
defparam \portB~16 .lut_mask = 16'hFF10;
defparam \portB~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N28
cycloneive_lcell_comb \portB~17 (
// Equation(s):
// \portB~17_combout  = (\portB~16_combout ) # ((dcifimemload_20 & (!cuifALUOP_21 & Mux391)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(\portB~16_combout ),
	.datad(Mux391),
	.cin(gnd),
	.combout(\portB~17_combout ),
	.cout());
// synopsys translate_off
defparam \portB~17 .lut_mask = 16'hF2F0;
defparam \portB~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N24
cycloneive_lcell_comb \portB~18 (
// Equation(s):
// \portB~18_combout  = (\portB~1_combout ) # ((!dcifimemload_20 & (!cuifALUOP_21 & Mux40)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux40),
	.datad(\portB~1_combout ),
	.cin(gnd),
	.combout(\portB~18_combout ),
	.cout());
// synopsys translate_off
defparam \portB~18 .lut_mask = 16'hFF10;
defparam \portB~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N16
cycloneive_lcell_comb \portB~19 (
// Equation(s):
// \portB~19_combout  = (\portB~18_combout ) # ((dcifimemload_20 & (!cuifALUOP_21 & Mux401)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux401),
	.datad(\portB~18_combout ),
	.cin(gnd),
	.combout(\portB~19_combout ),
	.cout());
// synopsys translate_off
defparam \portB~19 .lut_mask = 16'hFF20;
defparam \portB~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N20
cycloneive_lcell_comb \portB~20 (
// Equation(s):
// \portB~20_combout  = (\portB~1_combout ) # ((!cuifALUOP_21 & (!dcifimemload_20 & Mux41)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(Mux41),
	.datad(\portB~1_combout ),
	.cin(gnd),
	.combout(\portB~20_combout ),
	.cout());
// synopsys translate_off
defparam \portB~20 .lut_mask = 16'hFF10;
defparam \portB~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N18
cycloneive_lcell_comb \portB~21 (
// Equation(s):
// \portB~21_combout  = (\portB~20_combout ) # ((!cuifALUOP_21 & (Mux411 & dcifimemload_20)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(Mux411),
	.datac(dcifimemload_20),
	.datad(\portB~20_combout ),
	.cin(gnd),
	.combout(\portB~21_combout ),
	.cout());
// synopsys translate_off
defparam \portB~21 .lut_mask = 16'hFF40;
defparam \portB~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N20
cycloneive_lcell_comb \portB~22 (
// Equation(s):
// \portB~22_combout  = (\portB~1_combout ) # ((!cuifALUOP_21 & (!dcifimemload_20 & Mux42)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(\portB~1_combout ),
	.datad(Mux42),
	.cin(gnd),
	.combout(\portB~22_combout ),
	.cout());
// synopsys translate_off
defparam \portB~22 .lut_mask = 16'hF1F0;
defparam \portB~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N26
cycloneive_lcell_comb \portB~23 (
// Equation(s):
// \portB~23_combout  = (\portB~22_combout ) # ((!cuifALUOP_21 & (dcifimemload_20 & Mux421)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(Mux421),
	.datad(\portB~22_combout ),
	.cin(gnd),
	.combout(\portB~23_combout ),
	.cout());
// synopsys translate_off
defparam \portB~23 .lut_mask = 16'hFF40;
defparam \portB~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N24
cycloneive_lcell_comb \portB~24 (
// Equation(s):
// \portB~24_combout  = (\portB~1_combout ) # ((!dcifimemload_20 & (!cuifALUOP_21 & Mux43)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux43),
	.datad(\portB~1_combout ),
	.cin(gnd),
	.combout(\portB~24_combout ),
	.cout());
// synopsys translate_off
defparam \portB~24 .lut_mask = 16'hFF10;
defparam \portB~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N18
cycloneive_lcell_comb \portB~25 (
// Equation(s):
// \portB~25_combout  = (\portB~24_combout ) # ((!cuifALUOP_21 & (Mux431 & dcifimemload_20)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(Mux431),
	.datac(dcifimemload_20),
	.datad(\portB~24_combout ),
	.cin(gnd),
	.combout(\portB~25_combout ),
	.cout());
// synopsys translate_off
defparam \portB~25 .lut_mask = 16'hFF40;
defparam \portB~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N16
cycloneive_lcell_comb \portB~26 (
// Equation(s):
// \portB~26_combout  = (\portB~1_combout ) # ((!dcifimemload_20 & (!cuifALUOP_21 & Mux44)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux44),
	.datad(\portB~1_combout ),
	.cin(gnd),
	.combout(\portB~26_combout ),
	.cout());
// synopsys translate_off
defparam \portB~26 .lut_mask = 16'hFF10;
defparam \portB~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N14
cycloneive_lcell_comb \portB~27 (
// Equation(s):
// \portB~27_combout  = (\portB~26_combout ) # ((dcifimemload_20 & (Mux441 & !cuifALUOP_21)))

	.dataa(dcifimemload_20),
	.datab(Mux441),
	.datac(\CU|cuif.ALUOP[2]~20_combout ),
	.datad(\portB~26_combout ),
	.cin(gnd),
	.combout(\portB~27_combout ),
	.cout());
// synopsys translate_off
defparam \portB~27 .lut_mask = 16'hFF08;
defparam \portB~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N16
cycloneive_lcell_comb \portB~28 (
// Equation(s):
// \portB~28_combout  = (\portB~1_combout ) # ((!dcifimemload_20 & (!cuifALUOP_21 & Mux45)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux45),
	.datad(\portB~1_combout ),
	.cin(gnd),
	.combout(\portB~28_combout ),
	.cout());
// synopsys translate_off
defparam \portB~28 .lut_mask = 16'hFF10;
defparam \portB~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N30
cycloneive_lcell_comb \portB~29 (
// Equation(s):
// \portB~29_combout  = (\portB~28_combout ) # ((dcifimemload_20 & (!cuifALUOP_21 & Mux451)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux451),
	.datad(\portB~28_combout ),
	.cin(gnd),
	.combout(\portB~29_combout ),
	.cout());
// synopsys translate_off
defparam \portB~29 .lut_mask = 16'hFF20;
defparam \portB~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N2
cycloneive_lcell_comb \portB~30 (
// Equation(s):
// \portB~30_combout  = (\portB~1_combout ) # ((!cuifALUOP_21 & (!dcifimemload_20 & Mux46)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(\portB~1_combout ),
	.datad(Mux46),
	.cin(gnd),
	.combout(\portB~30_combout ),
	.cout());
// synopsys translate_off
defparam \portB~30 .lut_mask = 16'hF1F0;
defparam \portB~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N16
cycloneive_lcell_comb \portB~31 (
// Equation(s):
// \portB~31_combout  = (\portB~30_combout ) # ((!cuifALUOP_21 & (dcifimemload_20 & Mux461)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(Mux461),
	.datad(\portB~30_combout ),
	.cin(gnd),
	.combout(\portB~31_combout ),
	.cout());
// synopsys translate_off
defparam \portB~31 .lut_mask = 16'hFF40;
defparam \portB~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N6
cycloneive_lcell_comb \portB~32 (
// Equation(s):
// \portB~32_combout  = (\portB~1_combout ) # ((!cuifALUOP_21 & (!dcifimemload_20 & Mux47)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(\portB~1_combout ),
	.datad(Mux47),
	.cin(gnd),
	.combout(\portB~32_combout ),
	.cout());
// synopsys translate_off
defparam \portB~32 .lut_mask = 16'hF1F0;
defparam \portB~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N0
cycloneive_lcell_comb \portB~33 (
// Equation(s):
// \portB~33_combout  = (\portB~32_combout ) # ((!cuifALUOP_21 & (dcifimemload_20 & Mux471)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(Mux471),
	.datad(\portB~32_combout ),
	.cin(gnd),
	.combout(\portB~33_combout ),
	.cout());
// synopsys translate_off
defparam \portB~33 .lut_mask = 16'hFF40;
defparam \portB~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N18
cycloneive_lcell_comb \portB~34 (
// Equation(s):
// \portB~34_combout  = (\portB~0_combout ) # ((!cuifALUOP_21 & (!dcifimemload_20 & Mux48)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(\portB~0_combout ),
	.datad(Mux48),
	.cin(gnd),
	.combout(\portB~34_combout ),
	.cout());
// synopsys translate_off
defparam \portB~34 .lut_mask = 16'hF1F0;
defparam \portB~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N2
cycloneive_lcell_comb \portB~35 (
// Equation(s):
// \portB~35_combout  = (\portB~34_combout ) # ((!cuifALUOP_21 & (dcifimemload_20 & Mux481)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(Mux481),
	.datad(\portB~34_combout ),
	.cin(gnd),
	.combout(\portB~35_combout ),
	.cout());
// synopsys translate_off
defparam \portB~35 .lut_mask = 16'hFF40;
defparam \portB~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N6
cycloneive_lcell_comb \portB~36 (
// Equation(s):
// \portB~36_combout  = (cuifALUOP_21 & (((dcifimemload_14)))) # (!cuifALUOP_21 & (!dcifimemload_20 & ((Mux49))))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(dcifimemload_14),
	.datad(Mux49),
	.cin(gnd),
	.combout(\portB~36_combout ),
	.cout());
// synopsys translate_off
defparam \portB~36 .lut_mask = 16'hD1C0;
defparam \portB~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N30
cycloneive_lcell_comb \portB~37 (
// Equation(s):
// \portB~37_combout  = (\portB~36_combout ) # ((dcifimemload_20 & (!cuifALUOP_21 & Mux491)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux491),
	.datad(\portB~36_combout ),
	.cin(gnd),
	.combout(\portB~37_combout ),
	.cout());
// synopsys translate_off
defparam \portB~37 .lut_mask = 16'hFF20;
defparam \portB~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N10
cycloneive_lcell_comb \portB~38 (
// Equation(s):
// \portB~38_combout  = (cuifALUOP_21 & (dcifimemload_13)) # (!cuifALUOP_21 & (((!dcifimemload_20 & Mux50))))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_13),
	.datac(dcifimemload_20),
	.datad(Mux50),
	.cin(gnd),
	.combout(\portB~38_combout ),
	.cout());
// synopsys translate_off
defparam \portB~38 .lut_mask = 16'h8D88;
defparam \portB~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N20
cycloneive_lcell_comb \portB~39 (
// Equation(s):
// \portB~39_combout  = (\portB~38_combout ) # ((!cuifALUOP_21 & (dcifimemload_20 & Mux501)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(Mux501),
	.datad(\portB~38_combout ),
	.cin(gnd),
	.combout(\portB~39_combout ),
	.cout());
// synopsys translate_off
defparam \portB~39 .lut_mask = 16'hFF40;
defparam \portB~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N4
cycloneive_lcell_comb \portB~40 (
// Equation(s):
// \portB~40_combout  = (cuifALUOP_21 & (((dcifimemload_12)))) # (!cuifALUOP_21 & (!dcifimemload_20 & ((Mux51))))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(dcifimemload_12),
	.datad(Mux51),
	.cin(gnd),
	.combout(\portB~40_combout ),
	.cout());
// synopsys translate_off
defparam \portB~40 .lut_mask = 16'hB1A0;
defparam \portB~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N8
cycloneive_lcell_comb \portB~41 (
// Equation(s):
// \portB~41_combout  = (\portB~40_combout ) # ((!cuifALUOP_21 & (dcifimemload_20 & Mux511)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(\portB~40_combout ),
	.datad(Mux511),
	.cin(gnd),
	.combout(\portB~41_combout ),
	.cout());
// synopsys translate_off
defparam \portB~41 .lut_mask = 16'hF4F0;
defparam \portB~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N4
cycloneive_lcell_comb \portB~42 (
// Equation(s):
// \portB~42_combout  = (cuifALUOP_21 & (((dcifimemload_11)))) # (!cuifALUOP_21 & (!dcifimemload_20 & ((Mux52))))

	.dataa(dcifimemload_20),
	.datab(dcifimemload_11),
	.datac(\CU|cuif.ALUOP[2]~20_combout ),
	.datad(Mux52),
	.cin(gnd),
	.combout(\portB~42_combout ),
	.cout());
// synopsys translate_off
defparam \portB~42 .lut_mask = 16'hC5C0;
defparam \portB~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N6
cycloneive_lcell_comb \portB~43 (
// Equation(s):
// \portB~43_combout  = (\portB~42_combout ) # ((!cuifALUOP_21 & (dcifimemload_20 & Mux521)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(\portB~42_combout ),
	.datad(Mux521),
	.cin(gnd),
	.combout(\portB~43_combout ),
	.cout());
// synopsys translate_off
defparam \portB~43 .lut_mask = 16'hF4F0;
defparam \portB~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N30
cycloneive_lcell_comb \portB~44 (
// Equation(s):
// \portB~44_combout  = (cuifALUOP_21 & (((dcifimemload_10)))) # (!cuifALUOP_21 & (!dcifimemload_20 & ((Mux53))))

	.dataa(dcifimemload_20),
	.datab(dcifimemload_10),
	.datac(\CU|cuif.ALUOP[2]~20_combout ),
	.datad(Mux53),
	.cin(gnd),
	.combout(\portB~44_combout ),
	.cout());
// synopsys translate_off
defparam \portB~44 .lut_mask = 16'hC5C0;
defparam \portB~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N16
cycloneive_lcell_comb \portB~45 (
// Equation(s):
// \portB~45_combout  = (\portB~44_combout ) # ((!cuifALUOP_21 & (dcifimemload_20 & Mux531)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(\portB~44_combout ),
	.datad(Mux531),
	.cin(gnd),
	.combout(\portB~45_combout ),
	.cout());
// synopsys translate_off
defparam \portB~45 .lut_mask = 16'hF4F0;
defparam \portB~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N22
cycloneive_lcell_comb \portB~46 (
// Equation(s):
// \portB~46_combout  = (cuifALUOP_21 & (((dcifimemload_9)))) # (!cuifALUOP_21 & (!dcifimemload_20 & ((Mux54))))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(dcifimemload_9),
	.datad(Mux54),
	.cin(gnd),
	.combout(\portB~46_combout ),
	.cout());
// synopsys translate_off
defparam \portB~46 .lut_mask = 16'hD1C0;
defparam \portB~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N4
cycloneive_lcell_comb \portB~47 (
// Equation(s):
// \portB~47_combout  = (\portB~46_combout ) # ((dcifimemload_20 & (!cuifALUOP_21 & Mux541)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(\portB~46_combout ),
	.datad(Mux541),
	.cin(gnd),
	.combout(\portB~47_combout ),
	.cout());
// synopsys translate_off
defparam \portB~47 .lut_mask = 16'hF2F0;
defparam \portB~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N26
cycloneive_lcell_comb \portB~48 (
// Equation(s):
// \portB~48_combout  = (cuifALUOP_21 & (dcifimemload_8)) # (!cuifALUOP_21 & (((!dcifimemload_20 & Mux55))))

	.dataa(dcifimemload_8),
	.datab(dcifimemload_20),
	.datac(\CU|cuif.ALUOP[2]~20_combout ),
	.datad(Mux55),
	.cin(gnd),
	.combout(\portB~48_combout ),
	.cout());
// synopsys translate_off
defparam \portB~48 .lut_mask = 16'hA3A0;
defparam \portB~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N24
cycloneive_lcell_comb \portB~49 (
// Equation(s):
// \portB~49_combout  = (\portB~48_combout ) # ((dcifimemload_20 & (!cuifALUOP_21 & Mux551)))

	.dataa(\portB~48_combout ),
	.datab(dcifimemload_20),
	.datac(\CU|cuif.ALUOP[2]~20_combout ),
	.datad(Mux551),
	.cin(gnd),
	.combout(\portB~49_combout ),
	.cout());
// synopsys translate_off
defparam \portB~49 .lut_mask = 16'hAEAA;
defparam \portB~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N18
cycloneive_lcell_comb \portB~50 (
// Equation(s):
// \portB~50_combout  = (cuifALUOP_21 & (dcifimemload_7)) # (!cuifALUOP_21 & (((!dcifimemload_20 & Mux56))))

	.dataa(dcifimemload_7),
	.datab(dcifimemload_20),
	.datac(\CU|cuif.ALUOP[2]~20_combout ),
	.datad(Mux56),
	.cin(gnd),
	.combout(\portB~50_combout ),
	.cout());
// synopsys translate_off
defparam \portB~50 .lut_mask = 16'hA3A0;
defparam \portB~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N0
cycloneive_lcell_comb \portB~51 (
// Equation(s):
// \portB~51_combout  = (\portB~50_combout ) # ((Mux561 & (dcifimemload_20 & !cuifALUOP_21)))

	.dataa(Mux561),
	.datab(dcifimemload_20),
	.datac(\CU|cuif.ALUOP[2]~20_combout ),
	.datad(\portB~50_combout ),
	.cin(gnd),
	.combout(\portB~51_combout ),
	.cout());
// synopsys translate_off
defparam \portB~51 .lut_mask = 16'hFF08;
defparam \portB~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N10
cycloneive_lcell_comb \portB~52 (
// Equation(s):
// \portB~52_combout  = (cuifALUOP_21 & (((dcifimemload_6)))) # (!cuifALUOP_21 & (!dcifimemload_20 & ((Mux57))))

	.dataa(dcifimemload_20),
	.datab(dcifimemload_6),
	.datac(\CU|cuif.ALUOP[2]~20_combout ),
	.datad(Mux57),
	.cin(gnd),
	.combout(\portB~52_combout ),
	.cout());
// synopsys translate_off
defparam \portB~52 .lut_mask = 16'hC5C0;
defparam \portB~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N12
cycloneive_lcell_comb \portB~53 (
// Equation(s):
// \portB~53_combout  = (\portB~52_combout ) # ((dcifimemload_20 & (!cuifALUOP_21 & Mux571)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux571),
	.datad(\portB~52_combout ),
	.cin(gnd),
	.combout(\portB~53_combout ),
	.cout());
// synopsys translate_off
defparam \portB~53 .lut_mask = 16'hFF20;
defparam \portB~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N24
cycloneive_lcell_comb \portB~54 (
// Equation(s):
// \portB~54_combout  = (cuifALUOP_21 & (((dcifimemload_5)))) # (!cuifALUOP_21 & (!dcifimemload_20 & ((Mux58))))

	.dataa(dcifimemload_20),
	.datab(dcifimemload_5),
	.datac(\CU|cuif.ALUOP[2]~20_combout ),
	.datad(Mux58),
	.cin(gnd),
	.combout(\portB~54_combout ),
	.cout());
// synopsys translate_off
defparam \portB~54 .lut_mask = 16'hC5C0;
defparam \portB~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N10
cycloneive_lcell_comb \portB~55 (
// Equation(s):
// \portB~55_combout  = (\portB~54_combout ) # ((dcifimemload_20 & (!cuifALUOP_21 & Mux581)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux581),
	.datad(\portB~54_combout ),
	.cin(gnd),
	.combout(\portB~55_combout ),
	.cout());
// synopsys translate_off
defparam \portB~55 .lut_mask = 16'hFF20;
defparam \portB~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N12
cycloneive_lcell_comb \portB~56 (
// Equation(s):
// \portB~56_combout  = (cuifALUOP_21 & (((dcifimemload_4)))) # (!cuifALUOP_21 & (!dcifimemload_20 & ((Mux59))))

	.dataa(dcifimemload_20),
	.datab(dcifimemload_4),
	.datac(\CU|cuif.ALUOP[2]~20_combout ),
	.datad(Mux59),
	.cin(gnd),
	.combout(\portB~56_combout ),
	.cout());
// synopsys translate_off
defparam \portB~56 .lut_mask = 16'hC5C0;
defparam \portB~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N30
cycloneive_lcell_comb \portB~57 (
// Equation(s):
// \portB~57_combout  = (\portB~56_combout ) # ((dcifimemload_20 & (!cuifALUOP_21 & Mux591)))

	.dataa(dcifimemload_20),
	.datab(\CU|cuif.ALUOP[2]~20_combout ),
	.datac(Mux591),
	.datad(\portB~56_combout ),
	.cin(gnd),
	.combout(\portB~57_combout ),
	.cout());
// synopsys translate_off
defparam \portB~57 .lut_mask = 16'hFF20;
defparam \portB~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N4
cycloneive_lcell_comb \portB~58 (
// Equation(s):
// \portB~58_combout  = (cuifALUOP_21 & ((dcifimemload_3))) # (!cuifALUOP_21 & (dcifimemload_20))

	.dataa(dcifimemload_20),
	.datab(gnd),
	.datac(dcifimemload_3),
	.datad(\CU|cuif.ALUOP[2]~20_combout ),
	.cin(gnd),
	.combout(\portB~58_combout ),
	.cout());
// synopsys translate_off
defparam \portB~58 .lut_mask = 16'hF0AA;
defparam \portB~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N22
cycloneive_lcell_comb \portB~59 (
// Equation(s):
// \portB~59_combout  = (cuifALUOP_21 & (\portB~58_combout )) # (!cuifALUOP_21 & ((\portB~58_combout  & ((Mux60))) # (!\portB~58_combout  & (Mux601))))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(\portB~58_combout ),
	.datac(Mux601),
	.datad(Mux60),
	.cin(gnd),
	.combout(\portB~59_combout ),
	.cout());
// synopsys translate_off
defparam \portB~59 .lut_mask = 16'hDC98;
defparam \portB~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N6
cycloneive_lcell_comb \portB~60 (
// Equation(s):
// \portB~60_combout  = (cuifALUOP_21 & (dcifimemload_2)) # (!cuifALUOP_21 & (((!dcifimemload_20 & Mux61))))

	.dataa(dcifimemload_2),
	.datab(dcifimemload_20),
	.datac(\CU|cuif.ALUOP[2]~20_combout ),
	.datad(Mux61),
	.cin(gnd),
	.combout(\portB~60_combout ),
	.cout());
// synopsys translate_off
defparam \portB~60 .lut_mask = 16'hA3A0;
defparam \portB~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N0
cycloneive_lcell_comb \portB~61 (
// Equation(s):
// \portB~61_combout  = (\portB~60_combout ) # ((!cuifALUOP_21 & (dcifimemload_20 & Mux611)))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(dcifimemload_20),
	.datac(Mux611),
	.datad(\portB~60_combout ),
	.cin(gnd),
	.combout(\portB~61_combout ),
	.cout());
// synopsys translate_off
defparam \portB~61 .lut_mask = 16'hFF40;
defparam \portB~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N4
cycloneive_lcell_comb \portB~62 (
// Equation(s):
// \portB~62_combout  = (cuifALUOP_21 & (dcifimemload_1)) # (!cuifALUOP_21 & ((dcifimemload_20)))

	.dataa(gnd),
	.datab(dcifimemload_1),
	.datac(dcifimemload_20),
	.datad(\CU|cuif.ALUOP[2]~20_combout ),
	.cin(gnd),
	.combout(\portB~62_combout ),
	.cout());
// synopsys translate_off
defparam \portB~62 .lut_mask = 16'hCCF0;
defparam \portB~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N26
cycloneive_lcell_comb \portB~63 (
// Equation(s):
// \portB~63_combout  = (cuifALUOP_21 & (\portB~62_combout )) # (!cuifALUOP_21 & ((\portB~62_combout  & (Mux62)) # (!\portB~62_combout  & ((Mux621)))))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(\portB~62_combout ),
	.datac(Mux62),
	.datad(Mux621),
	.cin(gnd),
	.combout(\portB~63_combout ),
	.cout());
// synopsys translate_off
defparam \portB~63 .lut_mask = 16'hD9C8;
defparam \portB~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N8
cycloneive_lcell_comb \portB~64 (
// Equation(s):
// \portB~64_combout  = (cuifALUOP_21 & ((dcifimemload_0))) # (!cuifALUOP_21 & (dcifimemload_20))

	.dataa(dcifimemload_20),
	.datab(gnd),
	.datac(\CU|cuif.ALUOP[2]~20_combout ),
	.datad(dcifimemload_0),
	.cin(gnd),
	.combout(\portB~64_combout ),
	.cout());
// synopsys translate_off
defparam \portB~64 .lut_mask = 16'hFA0A;
defparam \portB~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N2
cycloneive_lcell_comb \portB~65 (
// Equation(s):
// \portB~65_combout  = (cuifALUOP_21 & (\portB~64_combout )) # (!cuifALUOP_21 & ((\portB~64_combout  & ((Mux63))) # (!\portB~64_combout  & (Mux631))))

	.dataa(\CU|cuif.ALUOP[2]~20_combout ),
	.datab(\portB~64_combout ),
	.datac(Mux631),
	.datad(Mux63),
	.cin(gnd),
	.combout(\portB~65_combout ),
	.cout());
// synopsys translate_off
defparam \portB~65 .lut_mask = 16'hDC98;
defparam \portB~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N24
cycloneive_lcell_comb \wdat~0 (
// Equation(s):
// \wdat~0_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & (PC_0)) # (!cuifMemtoReg_1 & ((ramiframload_0)))))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(\CU|cuif.MemtoReg[0]~0_combout ),
	.datac(PC_0),
	.datad(ramiframload_0),
	.cin(gnd),
	.combout(\wdat~0_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~0 .lut_mask = 16'hC480;
defparam \wdat~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N10
cycloneive_lcell_comb \wdat~1 (
// Equation(s):
// \wdat~1_combout  = (\wdat~0_combout ) # ((!cuifMemtoReg_1 & (Selector311 & !cuifMemtoReg_0)))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(\wdat~0_combout ),
	.datac(\ALU|Selector31~12_combout ),
	.datad(\CU|cuif.MemtoReg[0]~0_combout ),
	.cin(gnd),
	.combout(\wdat~1_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~1 .lut_mask = 16'hCCDC;
defparam \wdat~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N24
cycloneive_lcell_comb \wsel~0 (
// Equation(s):
// \wsel~0_combout  = (Equal31) # ((Equal0 & (dcifimemload_15)) # (!Equal0 & ((dcifimemload_20))))

	.dataa(dcifimemload_15),
	.datab(dcifimemload_20),
	.datac(\CU|Equal3~1_combout ),
	.datad(\CU|Equal0~2_combout ),
	.cin(gnd),
	.combout(\wsel~0_combout ),
	.cout());
// synopsys translate_off
defparam \wsel~0 .lut_mask = 16'hFAFC;
defparam \wsel~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N22
cycloneive_lcell_comb \wsel~1 (
// Equation(s):
// \wsel~1_combout  = (Equal31) # ((Equal0 & ((dcifimemload_14))) # (!Equal0 & (dcifimemload_19)))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_14),
	.datac(\CU|Equal3~1_combout ),
	.datad(\CU|Equal0~2_combout ),
	.cin(gnd),
	.combout(\wsel~1_combout ),
	.cout());
// synopsys translate_off
defparam \wsel~1 .lut_mask = 16'hFCFA;
defparam \wsel~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N0
cycloneive_lcell_comb \wsel~2 (
// Equation(s):
// \wsel~2_combout  = (Equal31) # ((Equal0 & ((dcifimemload_11))) # (!Equal0 & (dcifimemload_16)))

	.dataa(\CU|Equal3~1_combout ),
	.datab(dcifimemload_16),
	.datac(dcifimemload_11),
	.datad(\CU|Equal0~2_combout ),
	.cin(gnd),
	.combout(\wsel~2_combout ),
	.cout());
// synopsys translate_off
defparam \wsel~2 .lut_mask = 16'hFAEE;
defparam \wsel~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N30
cycloneive_lcell_comb \wsel~3 (
// Equation(s):
// \wsel~3_combout  = (Equal31) # ((Equal0 & ((dcifimemload_13))) # (!Equal0 & (dcifimemload_18)))

	.dataa(\CU|Equal3~1_combout ),
	.datab(dcifimemload_18),
	.datac(dcifimemload_13),
	.datad(\CU|Equal0~2_combout ),
	.cin(gnd),
	.combout(\wsel~3_combout ),
	.cout());
// synopsys translate_off
defparam \wsel~3 .lut_mask = 16'hFAEE;
defparam \wsel~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N4
cycloneive_lcell_comb \wsel~4 (
// Equation(s):
// \wsel~4_combout  = (Equal31) # ((Equal0 & ((dcifimemload_12))) # (!Equal0 & (dcifimemload_17)))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_12),
	.datac(\CU|Equal3~1_combout ),
	.datad(\CU|Equal0~2_combout ),
	.cin(gnd),
	.combout(\wsel~4_combout ),
	.cout());
// synopsys translate_off
defparam \wsel~4 .lut_mask = 16'hFCFA;
defparam \wsel~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N0
cycloneive_lcell_comb \wdat~2 (
// Equation(s):
// \wdat~2_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & (PC_1)) # (!cuifMemtoReg_1 & ((ramiframload_1)))))

	.dataa(PC_1),
	.datab(ramiframload_1),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(\CU|cuif.MemtoReg[1]~1_combout ),
	.cin(gnd),
	.combout(\wdat~2_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~2 .lut_mask = 16'hA0C0;
defparam \wdat~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N28
cycloneive_lcell_comb \wdat~3 (
// Equation(s):
// \wdat~3_combout  = (\wdat~2_combout ) # ((!cuifMemtoReg_0 & (!cuifMemtoReg_1 & Selector30)))

	.dataa(\CU|cuif.MemtoReg[0]~0_combout ),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\wdat~2_combout ),
	.datad(Selector30),
	.cin(gnd),
	.combout(\wdat~3_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~3 .lut_mask = 16'hF1F0;
defparam \wdat~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N20
cycloneive_lcell_comb \wdat~4 (
// Equation(s):
// \wdat~4_combout  = (cuifMemtoReg_1 & (cuifMemtoReg_0)) # (!cuifMemtoReg_1 & ((cuifMemtoReg_0 & (ramiframload_31)) # (!cuifMemtoReg_0 & ((Selector0)))))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(\CU|cuif.MemtoReg[0]~0_combout ),
	.datac(ramiframload_31),
	.datad(Selector0),
	.cin(gnd),
	.combout(\wdat~4_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~4 .lut_mask = 16'hD9C8;
defparam \wdat~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N22
cycloneive_lcell_comb \wdat~5 (
// Equation(s):
// \wdat~5_combout  = (cuifMemtoReg_1 & ((\wdat~4_combout  & ((\Add0~58_combout ))) # (!\wdat~4_combout  & (dcifimemload_15)))) # (!cuifMemtoReg_1 & (((\wdat~4_combout ))))

	.dataa(dcifimemload_15),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\Add0~58_combout ),
	.datad(\wdat~4_combout ),
	.cin(gnd),
	.combout(\wdat~5_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~5 .lut_mask = 16'hF388;
defparam \wdat~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N4
cycloneive_lcell_comb \wdat~6 (
// Equation(s):
// \wdat~6_combout  = (cuifMemtoReg_0 & ((ramiframload_30) # ((cuifMemtoReg_1)))) # (!cuifMemtoReg_0 & (((!cuifMemtoReg_1 & Selector1))))

	.dataa(\CU|cuif.MemtoReg[0]~0_combout ),
	.datab(ramiframload_30),
	.datac(\CU|cuif.MemtoReg[1]~1_combout ),
	.datad(Selector1),
	.cin(gnd),
	.combout(\wdat~6_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~6 .lut_mask = 16'hADA8;
defparam \wdat~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N6
cycloneive_lcell_comb \wdat~7 (
// Equation(s):
// \wdat~7_combout  = (cuifMemtoReg_1 & ((\wdat~6_combout  & (\Add0~56_combout )) # (!\wdat~6_combout  & ((dcifimemload_14))))) # (!cuifMemtoReg_1 & (((\wdat~6_combout ))))

	.dataa(\Add0~56_combout ),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\wdat~6_combout ),
	.datad(dcifimemload_14),
	.cin(gnd),
	.combout(\wdat~7_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~7 .lut_mask = 16'hBCB0;
defparam \wdat~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N18
cycloneive_lcell_comb \wdat~8 (
// Equation(s):
// \wdat~8_combout  = (cuifMemtoReg_1 & (cuifMemtoReg_0)) # (!cuifMemtoReg_1 & ((cuifMemtoReg_0 & (ramiframload_29)) # (!cuifMemtoReg_0 & ((Selector2)))))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(\CU|cuif.MemtoReg[0]~0_combout ),
	.datac(ramiframload_29),
	.datad(Selector2),
	.cin(gnd),
	.combout(\wdat~8_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~8 .lut_mask = 16'hD9C8;
defparam \wdat~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N20
cycloneive_lcell_comb \wdat~9 (
// Equation(s):
// \wdat~9_combout  = (cuifMemtoReg_1 & ((\wdat~8_combout  & (\Add0~54_combout )) # (!\wdat~8_combout  & ((dcifimemload_13))))) # (!cuifMemtoReg_1 & (((\wdat~8_combout ))))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(\Add0~54_combout ),
	.datac(dcifimemload_13),
	.datad(\wdat~8_combout ),
	.cin(gnd),
	.combout(\wdat~9_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~9 .lut_mask = 16'hDDA0;
defparam \wdat~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N14
cycloneive_lcell_comb \wdat~10 (
// Equation(s):
// \wdat~10_combout  = (cuifMemtoReg_1 & (((cuifMemtoReg_0)))) # (!cuifMemtoReg_1 & ((cuifMemtoReg_0 & (ramiframload_28)) # (!cuifMemtoReg_0 & ((Selector3)))))

	.dataa(ramiframload_28),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\wdat~10_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~10 .lut_mask = 16'hE3E0;
defparam \wdat~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N12
cycloneive_lcell_comb \wdat~11 (
// Equation(s):
// \wdat~11_combout  = (\wdat~10_combout  & ((\Add0~52_combout ) # ((!cuifMemtoReg_1)))) # (!\wdat~10_combout  & (((dcifimemload_12 & cuifMemtoReg_1))))

	.dataa(\Add0~52_combout ),
	.datab(dcifimemload_12),
	.datac(\wdat~10_combout ),
	.datad(\CU|cuif.MemtoReg[1]~1_combout ),
	.cin(gnd),
	.combout(\wdat~11_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~11 .lut_mask = 16'hACF0;
defparam \wdat~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N6
cycloneive_lcell_comb \wdat~12 (
// Equation(s):
// \wdat~12_combout  = (cuifMemtoReg_1 & (((cuifMemtoReg_0)))) # (!cuifMemtoReg_1 & ((cuifMemtoReg_0 & (ramiframload_27)) # (!cuifMemtoReg_0 & ((Selector41)))))

	.dataa(ramiframload_27),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\wdat~12_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~12 .lut_mask = 16'hE3E0;
defparam \wdat~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N24
cycloneive_lcell_comb \wdat~13 (
// Equation(s):
// \wdat~13_combout  = (cuifMemtoReg_1 & ((\wdat~12_combout  & ((\Add0~50_combout ))) # (!\wdat~12_combout  & (dcifimemload_11)))) # (!cuifMemtoReg_1 & (((\wdat~12_combout ))))

	.dataa(dcifimemload_11),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\Add0~50_combout ),
	.datad(\wdat~12_combout ),
	.cin(gnd),
	.combout(\wdat~13_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~13 .lut_mask = 16'hF388;
defparam \wdat~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N18
cycloneive_lcell_comb \wdat~14 (
// Equation(s):
// \wdat~14_combout  = (cuifMemtoReg_1 & (((cuifMemtoReg_0)))) # (!cuifMemtoReg_1 & ((cuifMemtoReg_0 & (ramiframload_26)) # (!cuifMemtoReg_0 & ((Selector51)))))

	.dataa(ramiframload_26),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(\ALU|Selector5~8_combout ),
	.cin(gnd),
	.combout(\wdat~14_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~14 .lut_mask = 16'hE3E0;
defparam \wdat~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N10
cycloneive_lcell_comb \wdat~15 (
// Equation(s):
// \wdat~15_combout  = (cuifMemtoReg_1 & ((\wdat~14_combout  & ((\Add0~48_combout ))) # (!\wdat~14_combout  & (dcifimemload_10)))) # (!cuifMemtoReg_1 & (((\wdat~14_combout ))))

	.dataa(dcifimemload_10),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\Add0~48_combout ),
	.datad(\wdat~14_combout ),
	.cin(gnd),
	.combout(\wdat~15_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~15 .lut_mask = 16'hF388;
defparam \wdat~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N10
cycloneive_lcell_comb \wdat~16 (
// Equation(s):
// \wdat~16_combout  = (cuifMemtoReg_1 & (((cuifMemtoReg_0)))) # (!cuifMemtoReg_1 & ((cuifMemtoReg_0 & (ramiframload_25)) # (!cuifMemtoReg_0 & ((Selector6)))))

	.dataa(ramiframload_25),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(Selector6),
	.datad(\CU|cuif.MemtoReg[0]~0_combout ),
	.cin(gnd),
	.combout(\wdat~16_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~16 .lut_mask = 16'hEE30;
defparam \wdat~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N16
cycloneive_lcell_comb \wdat~17 (
// Equation(s):
// \wdat~17_combout  = (cuifMemtoReg_1 & ((\wdat~16_combout  & (\Add0~46_combout )) # (!\wdat~16_combout  & ((dcifimemload_9))))) # (!cuifMemtoReg_1 & (((\wdat~16_combout ))))

	.dataa(\Add0~46_combout ),
	.datab(dcifimemload_9),
	.datac(\CU|cuif.MemtoReg[1]~1_combout ),
	.datad(\wdat~16_combout ),
	.cin(gnd),
	.combout(\wdat~17_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~17 .lut_mask = 16'hAFC0;
defparam \wdat~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N8
cycloneive_lcell_comb \wdat~18 (
// Equation(s):
// \wdat~18_combout  = (cuifMemtoReg_0 & ((ramiframload_24) # ((cuifMemtoReg_1)))) # (!cuifMemtoReg_0 & (((!cuifMemtoReg_1 & Selector7))))

	.dataa(\CU|cuif.MemtoReg[0]~0_combout ),
	.datab(ramiframload_24),
	.datac(\CU|cuif.MemtoReg[1]~1_combout ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\wdat~18_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~18 .lut_mask = 16'hADA8;
defparam \wdat~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N0
cycloneive_lcell_comb \wdat~19 (
// Equation(s):
// \wdat~19_combout  = (\wdat~18_combout  & ((\Add0~44_combout ) # ((!cuifMemtoReg_1)))) # (!\wdat~18_combout  & (((dcifimemload_8 & cuifMemtoReg_1))))

	.dataa(\Add0~44_combout ),
	.datab(dcifimemload_8),
	.datac(\wdat~18_combout ),
	.datad(\CU|cuif.MemtoReg[1]~1_combout ),
	.cin(gnd),
	.combout(\wdat~19_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~19 .lut_mask = 16'hACF0;
defparam \wdat~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N6
cycloneive_lcell_comb \wdat~20 (
// Equation(s):
// \wdat~20_combout  = (cuifMemtoReg_0 & ((ramiframload_23) # ((cuifMemtoReg_1)))) # (!cuifMemtoReg_0 & (((!cuifMemtoReg_1 & Selector84))))

	.dataa(\CU|cuif.MemtoReg[0]~0_combout ),
	.datab(ramiframload_23),
	.datac(\CU|cuif.MemtoReg[1]~1_combout ),
	.datad(\ALU|Selector8~10_combout ),
	.cin(gnd),
	.combout(\wdat~20_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~20 .lut_mask = 16'hADA8;
defparam \wdat~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N30
cycloneive_lcell_comb \wdat~21 (
// Equation(s):
// \wdat~21_combout  = (cuifMemtoReg_1 & ((\wdat~20_combout  & ((\Add0~42_combout ))) # (!\wdat~20_combout  & (dcifimemload_7)))) # (!cuifMemtoReg_1 & (((\wdat~20_combout ))))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(dcifimemload_7),
	.datac(\Add0~42_combout ),
	.datad(\wdat~20_combout ),
	.cin(gnd),
	.combout(\wdat~21_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~21 .lut_mask = 16'hF588;
defparam \wdat~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N0
cycloneive_lcell_comb \wdat~22 (
// Equation(s):
// \wdat~22_combout  = (cuifMemtoReg_0 & ((ramiframload_22) # ((cuifMemtoReg_1)))) # (!cuifMemtoReg_0 & (((!cuifMemtoReg_1 & Selector93))))

	.dataa(\CU|cuif.MemtoReg[0]~0_combout ),
	.datab(ramiframload_22),
	.datac(\CU|cuif.MemtoReg[1]~1_combout ),
	.datad(\ALU|Selector9~8_combout ),
	.cin(gnd),
	.combout(\wdat~22_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~22 .lut_mask = 16'hADA8;
defparam \wdat~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N2
cycloneive_lcell_comb \wdat~23 (
// Equation(s):
// \wdat~23_combout  = (cuifMemtoReg_1 & ((\wdat~22_combout  & ((\Add0~40_combout ))) # (!\wdat~22_combout  & (dcifimemload_6)))) # (!cuifMemtoReg_1 & (((\wdat~22_combout ))))

	.dataa(dcifimemload_6),
	.datab(\Add0~40_combout ),
	.datac(\CU|cuif.MemtoReg[1]~1_combout ),
	.datad(\wdat~22_combout ),
	.cin(gnd),
	.combout(\wdat~23_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~23 .lut_mask = 16'hCFA0;
defparam \wdat~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N30
cycloneive_lcell_comb \wdat~24 (
// Equation(s):
// \wdat~24_combout  = (cuifMemtoReg_1 & (((cuifMemtoReg_0)))) # (!cuifMemtoReg_1 & ((cuifMemtoReg_0 & (ramiframload_21)) # (!cuifMemtoReg_0 & ((Selector103)))))

	.dataa(ramiframload_21),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(\ALU|Selector10~8_combout ),
	.cin(gnd),
	.combout(\wdat~24_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~24 .lut_mask = 16'hE3E0;
defparam \wdat~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N0
cycloneive_lcell_comb \wdat~25 (
// Equation(s):
// \wdat~25_combout  = (cuifMemtoReg_1 & ((\wdat~24_combout  & (\Add0~38_combout )) # (!\wdat~24_combout  & ((dcifimemload_5))))) # (!cuifMemtoReg_1 & (((\wdat~24_combout ))))

	.dataa(\Add0~38_combout ),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(dcifimemload_5),
	.datad(\wdat~24_combout ),
	.cin(gnd),
	.combout(\wdat~25_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~25 .lut_mask = 16'hBBC0;
defparam \wdat~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N20
cycloneive_lcell_comb \wdat~26 (
// Equation(s):
// \wdat~26_combout  = (cuifMemtoReg_1 & (((cuifMemtoReg_0)))) # (!cuifMemtoReg_1 & ((cuifMemtoReg_0 & (ramiframload_20)) # (!cuifMemtoReg_0 & ((Selector111)))))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(ramiframload_20),
	.datac(\ALU|Selector11~9_combout ),
	.datad(\CU|cuif.MemtoReg[0]~0_combout ),
	.cin(gnd),
	.combout(\wdat~26_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~26 .lut_mask = 16'hEE50;
defparam \wdat~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N2
cycloneive_lcell_comb \wdat~27 (
// Equation(s):
// \wdat~27_combout  = (cuifMemtoReg_1 & ((\wdat~26_combout  & (\Add0~36_combout )) # (!\wdat~26_combout  & ((dcifimemload_4))))) # (!cuifMemtoReg_1 & (((\wdat~26_combout ))))

	.dataa(\Add0~36_combout ),
	.datab(dcifimemload_4),
	.datac(\CU|cuif.MemtoReg[1]~1_combout ),
	.datad(\wdat~26_combout ),
	.cin(gnd),
	.combout(\wdat~27_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~27 .lut_mask = 16'hAFC0;
defparam \wdat~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N6
cycloneive_lcell_comb \wdat~28 (
// Equation(s):
// \wdat~28_combout  = (cuifMemtoReg_1 & (((cuifMemtoReg_0)))) # (!cuifMemtoReg_1 & ((cuifMemtoReg_0 & (ramiframload_19)) # (!cuifMemtoReg_0 & ((Selector12)))))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(ramiframload_19),
	.datac(Selector12),
	.datad(\CU|cuif.MemtoReg[0]~0_combout ),
	.cin(gnd),
	.combout(\wdat~28_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~28 .lut_mask = 16'hEE50;
defparam \wdat~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N24
cycloneive_lcell_comb \wdat~29 (
// Equation(s):
// \wdat~29_combout  = (cuifMemtoReg_1 & ((\wdat~28_combout  & ((\Add0~34_combout ))) # (!\wdat~28_combout  & (dcifimemload_3)))) # (!cuifMemtoReg_1 & (((\wdat~28_combout ))))

	.dataa(dcifimemload_3),
	.datab(\Add0~34_combout ),
	.datac(\CU|cuif.MemtoReg[1]~1_combout ),
	.datad(\wdat~28_combout ),
	.cin(gnd),
	.combout(\wdat~29_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~29 .lut_mask = 16'hCFA0;
defparam \wdat~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N18
cycloneive_lcell_comb \wdat~30 (
// Equation(s):
// \wdat~30_combout  = (cuifMemtoReg_0 & ((ramiframload_18) # ((cuifMemtoReg_1)))) # (!cuifMemtoReg_0 & (((Selector13 & !cuifMemtoReg_1))))

	.dataa(\CU|cuif.MemtoReg[0]~0_combout ),
	.datab(ramiframload_18),
	.datac(Selector13),
	.datad(\CU|cuif.MemtoReg[1]~1_combout ),
	.cin(gnd),
	.combout(\wdat~30_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~30 .lut_mask = 16'hAAD8;
defparam \wdat~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N16
cycloneive_lcell_comb \wdat~31 (
// Equation(s):
// \wdat~31_combout  = (cuifMemtoReg_1 & ((\wdat~30_combout  & ((\Add0~32_combout ))) # (!\wdat~30_combout  & (dcifimemload_2)))) # (!cuifMemtoReg_1 & (((\wdat~30_combout ))))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(dcifimemload_2),
	.datac(\Add0~32_combout ),
	.datad(\wdat~30_combout ),
	.cin(gnd),
	.combout(\wdat~31_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~31 .lut_mask = 16'hF588;
defparam \wdat~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N14
cycloneive_lcell_comb \wdat~32 (
// Equation(s):
// \wdat~32_combout  = (cuifMemtoReg_0 & ((ramiframload_17) # ((cuifMemtoReg_1)))) # (!cuifMemtoReg_0 & (((Selector143 & !cuifMemtoReg_1))))

	.dataa(\CU|cuif.MemtoReg[0]~0_combout ),
	.datab(ramiframload_17),
	.datac(\ALU|Selector14~8_combout ),
	.datad(\CU|cuif.MemtoReg[1]~1_combout ),
	.cin(gnd),
	.combout(\wdat~32_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~32 .lut_mask = 16'hAAD8;
defparam \wdat~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N12
cycloneive_lcell_comb \wdat~33 (
// Equation(s):
// \wdat~33_combout  = (\wdat~32_combout  & ((\Add0~30_combout ) # ((!cuifMemtoReg_1)))) # (!\wdat~32_combout  & (((dcifimemload_1 & cuifMemtoReg_1))))

	.dataa(\Add0~30_combout ),
	.datab(dcifimemload_1),
	.datac(\wdat~32_combout ),
	.datad(\CU|cuif.MemtoReg[1]~1_combout ),
	.cin(gnd),
	.combout(\wdat~33_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~33 .lut_mask = 16'hACF0;
defparam \wdat~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N30
cycloneive_lcell_comb \wdat~34 (
// Equation(s):
// \wdat~34_combout  = (cuifMemtoReg_1 & (cuifMemtoReg_0)) # (!cuifMemtoReg_1 & ((cuifMemtoReg_0 & (ramiframload_16)) # (!cuifMemtoReg_0 & ((Selector15)))))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(\CU|cuif.MemtoReg[0]~0_combout ),
	.datac(ramiframload_16),
	.datad(Selector15),
	.cin(gnd),
	.combout(\wdat~34_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~34 .lut_mask = 16'hD9C8;
defparam \wdat~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N26
cycloneive_lcell_comb \wdat~35 (
// Equation(s):
// \wdat~35_combout  = (\wdat~34_combout  & (((\Add0~28_combout ) # (!cuifMemtoReg_1)))) # (!\wdat~34_combout  & (dcifimemload_0 & (cuifMemtoReg_1)))

	.dataa(dcifimemload_0),
	.datab(\wdat~34_combout ),
	.datac(\CU|cuif.MemtoReg[1]~1_combout ),
	.datad(\Add0~28_combout ),
	.cin(gnd),
	.combout(\wdat~35_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~35 .lut_mask = 16'hEC2C;
defparam \wdat~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N18
cycloneive_lcell_comb \wdat~36 (
// Equation(s):
// \wdat~36_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & ((\Add0~26_combout ))) # (!cuifMemtoReg_1 & (ramiframload_15))))

	.dataa(ramiframload_15),
	.datab(\Add0~26_combout ),
	.datac(\CU|cuif.MemtoReg[1]~1_combout ),
	.datad(\CU|cuif.MemtoReg[0]~0_combout ),
	.cin(gnd),
	.combout(\wdat~36_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~36 .lut_mask = 16'hCA00;
defparam \wdat~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N14
cycloneive_lcell_comb \wdat~37 (
// Equation(s):
// \wdat~37_combout  = (\wdat~36_combout ) # ((!cuifMemtoReg_1 & (!cuifMemtoReg_0 & Selector16)))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(\CU|cuif.MemtoReg[0]~0_combout ),
	.datac(\wdat~36_combout ),
	.datad(Selector16),
	.cin(gnd),
	.combout(\wdat~37_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~37 .lut_mask = 16'hF1F0;
defparam \wdat~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N20
cycloneive_lcell_comb \wdat~38 (
// Equation(s):
// \wdat~38_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & (\Add0~24_combout )) # (!cuifMemtoReg_1 & ((ramiframload_14)))))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(\Add0~24_combout ),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(ramiframload_14),
	.cin(gnd),
	.combout(\wdat~38_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~38 .lut_mask = 16'hD080;
defparam \wdat~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N6
cycloneive_lcell_comb \wdat~39 (
// Equation(s):
// \wdat~39_combout  = (\wdat~38_combout ) # ((!cuifMemtoReg_1 & (!cuifMemtoReg_0 & Selector17)))

	.dataa(\wdat~38_combout ),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(Selector17),
	.cin(gnd),
	.combout(\wdat~39_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~39 .lut_mask = 16'hABAA;
defparam \wdat~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N4
cycloneive_lcell_comb \wdat~40 (
// Equation(s):
// \wdat~40_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & (\Add0~22_combout )) # (!cuifMemtoReg_1 & ((ramiframload_13)))))

	.dataa(\Add0~22_combout ),
	.datab(\CU|cuif.MemtoReg[0]~0_combout ),
	.datac(ramiframload_13),
	.datad(\CU|cuif.MemtoReg[1]~1_combout ),
	.cin(gnd),
	.combout(\wdat~40_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~40 .lut_mask = 16'h88C0;
defparam \wdat~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N18
cycloneive_lcell_comb \wdat~41 (
// Equation(s):
// \wdat~41_combout  = (\wdat~40_combout ) # ((!cuifMemtoReg_1 & (!cuifMemtoReg_0 & Selector18)))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(\CU|cuif.MemtoReg[0]~0_combout ),
	.datac(\wdat~40_combout ),
	.datad(Selector18),
	.cin(gnd),
	.combout(\wdat~41_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~41 .lut_mask = 16'hF1F0;
defparam \wdat~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N28
cycloneive_lcell_comb \wdat~42 (
// Equation(s):
// \wdat~42_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & (\Add0~20_combout )) # (!cuifMemtoReg_1 & ((ramiframload_12)))))

	.dataa(\CU|cuif.MemtoReg[0]~0_combout ),
	.datab(\Add0~20_combout ),
	.datac(ramiframload_12),
	.datad(\CU|cuif.MemtoReg[1]~1_combout ),
	.cin(gnd),
	.combout(\wdat~42_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~42 .lut_mask = 16'h88A0;
defparam \wdat~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N22
cycloneive_lcell_comb \wdat~43 (
// Equation(s):
// \wdat~43_combout  = (\wdat~42_combout ) # ((!cuifMemtoReg_1 & (!cuifMemtoReg_0 & Selector19)))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(\CU|cuif.MemtoReg[0]~0_combout ),
	.datac(\wdat~42_combout ),
	.datad(Selector19),
	.cin(gnd),
	.combout(\wdat~43_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~43 .lut_mask = 16'hF1F0;
defparam \wdat~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N6
cycloneive_lcell_comb \wdat~44 (
// Equation(s):
// \wdat~44_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & (\Add0~18_combout )) # (!cuifMemtoReg_1 & ((ramiframload_11)))))

	.dataa(\Add0~18_combout ),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(ramiframload_11),
	.cin(gnd),
	.combout(\wdat~44_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~44 .lut_mask = 16'hB080;
defparam \wdat~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N4
cycloneive_lcell_comb \wdat~45 (
// Equation(s):
// \wdat~45_combout  = (\wdat~44_combout ) # ((!cuifMemtoReg_1 & (!cuifMemtoReg_0 & Selector203)))

	.dataa(\wdat~44_combout ),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(\ALU|Selector20~9_combout ),
	.cin(gnd),
	.combout(\wdat~45_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~45 .lut_mask = 16'hABAA;
defparam \wdat~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N22
cycloneive_lcell_comb \wdat~46 (
// Equation(s):
// \wdat~46_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & ((\Add0~16_combout ))) # (!cuifMemtoReg_1 & (ramiframload_10))))

	.dataa(ramiframload_10),
	.datab(\CU|cuif.MemtoReg[0]~0_combout ),
	.datac(\Add0~16_combout ),
	.datad(\CU|cuif.MemtoReg[1]~1_combout ),
	.cin(gnd),
	.combout(\wdat~46_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~46 .lut_mask = 16'hC088;
defparam \wdat~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N14
cycloneive_lcell_comb \wdat~47 (
// Equation(s):
// \wdat~47_combout  = (\wdat~46_combout ) # ((!cuifMemtoReg_0 & (!cuifMemtoReg_1 & Selector213)))

	.dataa(\CU|cuif.MemtoReg[0]~0_combout ),
	.datab(\wdat~46_combout ),
	.datac(\CU|cuif.MemtoReg[1]~1_combout ),
	.datad(\ALU|Selector21~8_combout ),
	.cin(gnd),
	.combout(\wdat~47_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~47 .lut_mask = 16'hCDCC;
defparam \wdat~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N12
cycloneive_lcell_comb \wdat~48 (
// Equation(s):
// \wdat~48_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & (\Add0~14_combout )) # (!cuifMemtoReg_1 & ((ramiframload_9)))))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(\Add0~14_combout ),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(ramiframload_9),
	.cin(gnd),
	.combout(\wdat~48_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~48 .lut_mask = 16'hD080;
defparam \wdat~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N18
cycloneive_lcell_comb \wdat~49 (
// Equation(s):
// \wdat~49_combout  = (\wdat~48_combout ) # ((!cuifMemtoReg_1 & (!cuifMemtoReg_0 & Selector221)))

	.dataa(\wdat~48_combout ),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(Selector221),
	.cin(gnd),
	.combout(\wdat~49_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~49 .lut_mask = 16'hABAA;
defparam \wdat~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N16
cycloneive_lcell_comb \wdat~50 (
// Equation(s):
// \wdat~50_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & ((\Add0~12_combout ))) # (!cuifMemtoReg_1 & (ramiframload_8))))

	.dataa(\CU|cuif.MemtoReg[0]~0_combout ),
	.datab(ramiframload_8),
	.datac(\Add0~12_combout ),
	.datad(\CU|cuif.MemtoReg[1]~1_combout ),
	.cin(gnd),
	.combout(\wdat~50_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~50 .lut_mask = 16'hA088;
defparam \wdat~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N30
cycloneive_lcell_comb \wdat~51 (
// Equation(s):
// \wdat~51_combout  = (\wdat~50_combout ) # ((!cuifMemtoReg_0 & (!cuifMemtoReg_1 & Selector233)))

	.dataa(\CU|cuif.MemtoReg[0]~0_combout ),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\wdat~50_combout ),
	.datad(\ALU|Selector23~11_combout ),
	.cin(gnd),
	.combout(\wdat~51_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~51 .lut_mask = 16'hF1F0;
defparam \wdat~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N30
cycloneive_lcell_comb \wdat~52 (
// Equation(s):
// \wdat~52_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & (\Add0~10_combout )) # (!cuifMemtoReg_1 & ((ramiframload_7)))))

	.dataa(\Add0~10_combout ),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(ramiframload_7),
	.cin(gnd),
	.combout(\wdat~52_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~52 .lut_mask = 16'hB080;
defparam \wdat~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N28
cycloneive_lcell_comb \wdat~53 (
// Equation(s):
// \wdat~53_combout  = (\wdat~52_combout ) # ((!cuifMemtoReg_0 & (Selector242 & !cuifMemtoReg_1)))

	.dataa(\CU|cuif.MemtoReg[0]~0_combout ),
	.datab(Selector242),
	.datac(\CU|cuif.MemtoReg[1]~1_combout ),
	.datad(\wdat~52_combout ),
	.cin(gnd),
	.combout(\wdat~53_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~53 .lut_mask = 16'hFF04;
defparam \wdat~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N8
cycloneive_lcell_comb \wdat~54 (
// Equation(s):
// \wdat~54_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & (\Add0~8_combout )) # (!cuifMemtoReg_1 & ((ramiframload_6)))))

	.dataa(\Add0~8_combout ),
	.datab(ramiframload_6),
	.datac(\CU|cuif.MemtoReg[1]~1_combout ),
	.datad(\CU|cuif.MemtoReg[0]~0_combout ),
	.cin(gnd),
	.combout(\wdat~54_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~54 .lut_mask = 16'hAC00;
defparam \wdat~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N14
cycloneive_lcell_comb \wdat~55 (
// Equation(s):
// \wdat~55_combout  = (\wdat~54_combout ) # ((!cuifMemtoReg_1 & (!cuifMemtoReg_0 & Selector25)))

	.dataa(\wdat~54_combout ),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(Selector25),
	.cin(gnd),
	.combout(\wdat~55_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~55 .lut_mask = 16'hABAA;
defparam \wdat~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N8
cycloneive_lcell_comb \wdat~56 (
// Equation(s):
// \wdat~56_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & ((\Add0~6_combout ))) # (!cuifMemtoReg_1 & (ramiframload_5))))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(ramiframload_5),
	.datac(\Add0~6_combout ),
	.datad(\CU|cuif.MemtoReg[0]~0_combout ),
	.cin(gnd),
	.combout(\wdat~56_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~56 .lut_mask = 16'hE400;
defparam \wdat~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N12
cycloneive_lcell_comb \wdat~57 (
// Equation(s):
// \wdat~57_combout  = (\wdat~56_combout ) # ((!cuifMemtoReg_0 & (!cuifMemtoReg_1 & Selector261)))

	.dataa(\CU|cuif.MemtoReg[0]~0_combout ),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\wdat~56_combout ),
	.datad(\ALU|Selector26~8_combout ),
	.cin(gnd),
	.combout(\wdat~57_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~57 .lut_mask = 16'hF1F0;
defparam \wdat~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N30
cycloneive_lcell_comb \wdat~58 (
// Equation(s):
// \wdat~58_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & ((\Add0~4_combout ))) # (!cuifMemtoReg_1 & (ramiframload_4))))

	.dataa(\CU|cuif.MemtoReg[1]~1_combout ),
	.datab(ramiframload_4),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(\Add0~4_combout ),
	.cin(gnd),
	.combout(\wdat~58_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~58 .lut_mask = 16'hE040;
defparam \wdat~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N22
cycloneive_lcell_comb \wdat~59 (
// Equation(s):
// \wdat~59_combout  = (\wdat~58_combout ) # ((!cuifMemtoReg_1 & (!cuifMemtoReg_0 & Selector27)))

	.dataa(\wdat~58_combout ),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(Selector27),
	.cin(gnd),
	.combout(\wdat~59_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~59 .lut_mask = 16'hABAA;
defparam \wdat~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N22
cycloneive_lcell_comb \wdat~60 (
// Equation(s):
// \wdat~60_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & ((\Add0~2_combout ))) # (!cuifMemtoReg_1 & (ramiframload_3))))

	.dataa(\CU|cuif.MemtoReg[0]~0_combout ),
	.datab(ramiframload_3),
	.datac(\Add0~2_combout ),
	.datad(\CU|cuif.MemtoReg[1]~1_combout ),
	.cin(gnd),
	.combout(\wdat~60_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~60 .lut_mask = 16'hA088;
defparam \wdat~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N26
cycloneive_lcell_comb \wdat~61 (
// Equation(s):
// \wdat~61_combout  = (\wdat~60_combout ) # ((!cuifMemtoReg_1 & (!cuifMemtoReg_0 & Selector28)))

	.dataa(\wdat~60_combout ),
	.datab(\CU|cuif.MemtoReg[1]~1_combout ),
	.datac(\CU|cuif.MemtoReg[0]~0_combout ),
	.datad(Selector28),
	.cin(gnd),
	.combout(\wdat~61_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~61 .lut_mask = 16'hABAA;
defparam \wdat~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N26
cycloneive_lcell_comb \wdat~62 (
// Equation(s):
// \wdat~62_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & ((\Add0~0_combout ))) # (!cuifMemtoReg_1 & (ramiframload_2))))

	.dataa(ramiframload_2),
	.datab(\Add0~0_combout ),
	.datac(\CU|cuif.MemtoReg[1]~1_combout ),
	.datad(\CU|cuif.MemtoReg[0]~0_combout ),
	.cin(gnd),
	.combout(\wdat~62_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~62 .lut_mask = 16'hCA00;
defparam \wdat~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N4
cycloneive_lcell_comb \wdat~63 (
// Equation(s):
// \wdat~63_combout  = (\wdat~62_combout ) # ((!cuifMemtoReg_0 & (!cuifMemtoReg_1 & Selector291)))

	.dataa(\wdat~62_combout ),
	.datab(\CU|cuif.MemtoReg[0]~0_combout ),
	.datac(\CU|cuif.MemtoReg[1]~1_combout ),
	.datad(\ALU|Selector29~8_combout ),
	.cin(gnd),
	.combout(\wdat~63_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~63 .lut_mask = 16'hABAA;
defparam \wdat~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: DDIOOUTCELL_X60_Y0_N18
dffeas \dpif.halt (
	.clk(CLK),
	.d(\CU|Equal6~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dpifhalt),
	.prn(vcc));
// synopsys translate_off
defparam \dpif.halt .is_wysiwyg = "true";
defparam \dpif.halt .power_up = "low";
// synopsys translate_on

endmodule

module alu (
	Mux30,
	Mux301,
	dcifimemload_25,
	Mux302,
	cuifALUOP_3,
	cuifALUOP_2,
	cuifALUOP_1,
	cuifALUOP_0,
	Mux0,
	portB,
	Mux1,
	portB1,
	Mux2,
	portB2,
	Mux3,
	portB3,
	Mux4,
	portB4,
	Mux5,
	portB5,
	Mux6,
	portB6,
	Mux7,
	Mux71,
	Mux72,
	portB7,
	Mux8,
	portB8,
	Mux9,
	portB9,
	Mux10,
	portB10,
	Mux11,
	portB11,
	Mux12,
	portB12,
	Mux13,
	portB13,
	Mux14,
	portB14,
	Mux15,
	portB15,
	Mux16,
	portB16,
	Mux17,
	portB17,
	Mux18,
	portB18,
	Mux19,
	portB19,
	Mux20,
	portB20,
	Mux21,
	portB21,
	Mux22,
	portB22,
	Mux23,
	portB23,
	Mux24,
	Mux241,
	Mux242,
	portB24,
	Mux25,
	Mux251,
	Mux252,
	portB25,
	Mux26,
	portB26,
	Mux27,
	Mux271,
	Mux272,
	portB27,
	Mux28,
	portB28,
	Mux29,
	Mux291,
	Mux292,
	portB29,
	portB30,
	Mux31,
	Mux311,
	Mux312,
	portB31,
	Selector31,
	ShiftRight0,
	Selector24,
	Selector8,
	Selector0,
	Selector3,
	Selector4,
	Selector7,
	Selector11,
	ShiftRight01,
	Selector111,
	Selector15,
	Selector22,
	Selector28,
	Selector29,
	ShiftRight02,
	ShiftRight03,
	Selector291,
	ShiftLeft0,
	Selector10,
	Selector101,
	Selector102,
	Selector103,
	Selector2,
	Selector1,
	Selector41,
	Selector5,
	Selector51,
	Selector12,
	Selector241,
	Selector242,
	Selector13,
	Selector25,
	Selector14,
	Selector141,
	Selector142,
	Selector143,
	Selector27,
	Selector16,
	Selector18,
	Selector17,
	Selector6,
	Selector26,
	Selector261,
	Selector19,
	Selector20,
	Selector201,
	Selector202,
	Selector21,
	Selector211,
	Selector212,
	Selector213,
	Selector81,
	Selector82,
	Selector83,
	Selector84,
	Selector9,
	Selector91,
	Selector92,
	Selector93,
	Selector221,
	Selector30,
	Selector23,
	Selector231,
	Selector232,
	Equal0,
	Selector203,
	Selector311,
	Selector233,
	devpor,
	devclrn,
	devoe);
input 	Mux30;
input 	Mux301;
input 	dcifimemload_25;
input 	Mux302;
input 	cuifALUOP_3;
input 	cuifALUOP_2;
input 	cuifALUOP_1;
input 	cuifALUOP_0;
input 	Mux0;
input 	portB;
input 	Mux1;
input 	portB1;
input 	Mux2;
input 	portB2;
input 	Mux3;
input 	portB3;
input 	Mux4;
input 	portB4;
input 	Mux5;
input 	portB5;
input 	Mux6;
input 	portB6;
input 	Mux7;
input 	Mux71;
input 	Mux72;
input 	portB7;
input 	Mux8;
input 	portB8;
input 	Mux9;
input 	portB9;
input 	Mux10;
input 	portB10;
input 	Mux11;
input 	portB11;
input 	Mux12;
input 	portB12;
input 	Mux13;
input 	portB13;
input 	Mux14;
input 	portB14;
input 	Mux15;
input 	portB15;
input 	Mux16;
input 	portB16;
input 	Mux17;
input 	portB17;
input 	Mux18;
input 	portB18;
input 	Mux19;
input 	portB19;
input 	Mux20;
input 	portB20;
input 	Mux21;
input 	portB21;
input 	Mux22;
input 	portB22;
input 	Mux23;
input 	portB23;
input 	Mux24;
input 	Mux241;
input 	Mux242;
input 	portB24;
input 	Mux25;
input 	Mux251;
input 	Mux252;
input 	portB25;
input 	Mux26;
input 	portB26;
input 	Mux27;
input 	Mux271;
input 	Mux272;
input 	portB27;
input 	Mux28;
input 	portB28;
input 	Mux29;
input 	Mux291;
input 	Mux292;
input 	portB29;
input 	portB30;
input 	Mux31;
input 	Mux311;
input 	Mux312;
input 	portB31;
output 	Selector31;
output 	ShiftRight0;
output 	Selector24;
output 	Selector8;
output 	Selector0;
output 	Selector3;
output 	Selector4;
output 	Selector7;
output 	Selector11;
output 	ShiftRight01;
output 	Selector111;
output 	Selector15;
output 	Selector22;
output 	Selector28;
output 	Selector29;
output 	ShiftRight02;
output 	ShiftRight03;
output 	Selector291;
output 	ShiftLeft0;
output 	Selector10;
output 	Selector101;
output 	Selector102;
output 	Selector103;
output 	Selector2;
output 	Selector1;
output 	Selector41;
output 	Selector5;
output 	Selector51;
output 	Selector12;
output 	Selector241;
output 	Selector242;
output 	Selector13;
output 	Selector25;
output 	Selector14;
output 	Selector141;
output 	Selector142;
output 	Selector143;
output 	Selector27;
output 	Selector16;
output 	Selector18;
output 	Selector17;
output 	Selector6;
output 	Selector26;
output 	Selector261;
output 	Selector19;
output 	Selector20;
output 	Selector201;
output 	Selector202;
output 	Selector21;
output 	Selector211;
output 	Selector212;
output 	Selector213;
output 	Selector81;
output 	Selector82;
output 	Selector83;
output 	Selector84;
output 	Selector9;
output 	Selector91;
output 	Selector92;
output 	Selector93;
output 	Selector221;
output 	Selector30;
output 	Selector23;
output 	Selector231;
output 	Selector232;
output 	Equal0;
output 	Selector203;
output 	Selector311;
output 	Selector233;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~26_combout ;
wire \Add0~2_combout ;
wire \ShiftRight0~15_combout ;
wire \ShiftRight0~21_combout ;
wire \Selector0~19_combout ;
wire \ShiftLeft0~14_combout ;
wire \Selector0~24_combout ;
wire \ShiftLeft0~25_combout ;
wire \ShiftLeft0~36_combout ;
wire \Selector0~34_combout ;
wire \ShiftRight0~56_combout ;
wire \ShiftRight0~79_combout ;
wire \Selector12~3_combout ;
wire \Selector12~4_combout ;
wire \Selector12~5_combout ;
wire \ShiftRight0~101_combout ;
wire \Selector13~3_combout ;
wire \Selector13~4_combout ;
wire \Selector13~5_combout ;
wire \ShiftRight0~104_combout ;
wire \Selector27~2_combout ;
wire \Selector18~3_combout ;
wire \Selector18~4_combout ;
wire \Selector18~5_combout ;
wire \Selector17~3_combout ;
wire \Selector17~4_combout ;
wire \Selector17~5_combout ;
wire \Selector0~4_combout ;
wire \Selector0~5_combout ;
wire \Selector0~6_combout ;
wire \Selector31~4_combout ;
wire \Add1~0_combout ;
wire \Selector0~8_combout ;
wire \ShiftRight0~23_combout ;
wire \Selector0~9_combout ;
wire \ShiftRight0~20_combout ;
wire \ShiftRight0~14_combout ;
wire \ShiftRight0~17_combout ;
wire \ShiftRight0~16_combout ;
wire \ShiftRight0~18_combout ;
wire \ShiftRight0~19_combout ;
wire \ShiftRight0~22_combout ;
wire \Selector31~11_combout ;
wire \Selector31~6_combout ;
wire \Selector31~5_combout ;
wire \Selector31~7_combout ;
wire \Selector0~12_combout ;
wire \Add0~0_combout ;
wire \Selector0~11_combout ;
wire \Selector31~8_combout ;
wire \LessThan0~1_cout ;
wire \LessThan0~3_cout ;
wire \LessThan0~5_cout ;
wire \LessThan0~7_cout ;
wire \LessThan0~9_cout ;
wire \LessThan0~11_cout ;
wire \LessThan0~13_cout ;
wire \LessThan0~15_cout ;
wire \LessThan0~17_cout ;
wire \LessThan0~19_cout ;
wire \LessThan0~21_cout ;
wire \LessThan0~23_cout ;
wire \LessThan0~25_cout ;
wire \LessThan0~27_cout ;
wire \LessThan0~29_cout ;
wire \LessThan0~31_cout ;
wire \LessThan0~33_cout ;
wire \LessThan0~35_cout ;
wire \LessThan0~37_cout ;
wire \LessThan0~39_cout ;
wire \LessThan0~41_cout ;
wire \LessThan0~43_cout ;
wire \LessThan0~45_cout ;
wire \LessThan0~47_cout ;
wire \LessThan0~49_cout ;
wire \LessThan0~51_cout ;
wire \LessThan0~53_cout ;
wire \LessThan0~55_cout ;
wire \LessThan0~57_cout ;
wire \LessThan0~59_cout ;
wire \LessThan0~61_cout ;
wire \LessThan0~62_combout ;
wire \Selector31~9_combout ;
wire \LessThan1~1_cout ;
wire \LessThan1~3_cout ;
wire \LessThan1~5_cout ;
wire \LessThan1~7_cout ;
wire \LessThan1~9_cout ;
wire \LessThan1~11_cout ;
wire \LessThan1~13_cout ;
wire \LessThan1~15_cout ;
wire \LessThan1~17_cout ;
wire \LessThan1~19_cout ;
wire \LessThan1~21_cout ;
wire \LessThan1~23_cout ;
wire \LessThan1~25_cout ;
wire \LessThan1~27_cout ;
wire \LessThan1~29_cout ;
wire \LessThan1~31_cout ;
wire \LessThan1~33_cout ;
wire \LessThan1~35_cout ;
wire \LessThan1~37_cout ;
wire \LessThan1~39_cout ;
wire \LessThan1~41_cout ;
wire \LessThan1~43_cout ;
wire \LessThan1~45_cout ;
wire \LessThan1~47_cout ;
wire \LessThan1~49_cout ;
wire \LessThan1~51_cout ;
wire \LessThan1~53_cout ;
wire \LessThan1~55_cout ;
wire \LessThan1~57_cout ;
wire \LessThan1~59_cout ;
wire \LessThan1~61_cout ;
wire \LessThan1~62_combout ;
wire \ShiftRight0~37_combout ;
wire \ShiftRight0~38_combout ;
wire \ShiftRight0~39_combout ;
wire \ShiftRight0~40_combout ;
wire \ShiftRight0~42_combout ;
wire \ShiftRight0~43_combout ;
wire \ShiftRight0~123_combout ;
wire \ShiftRight0~44_combout ;
wire \ShiftRight0~45_combout ;
wire \ShiftRight0~46_combout ;
wire \ShiftRight0~47_combout ;
wire \ShiftRight0~48_combout ;
wire \ShiftRight0~49_combout ;
wire \ShiftRight0~35_combout ;
wire \ShiftRight0~31_combout ;
wire \ShiftRight0~32_combout ;
wire \ShiftRight0~33_combout ;
wire \Selector23~2_combout ;
wire \ShiftRight0~24_combout ;
wire \ShiftRight0~25_combout ;
wire \ShiftRight0~26_combout ;
wire \ShiftRight0~122_combout ;
wire \ShiftRight0~27_combout ;
wire \ShiftRight0~28_combout ;
wire \ShiftRight0~29_combout ;
wire \ShiftRight0~30_combout ;
wire \ShiftRight0~36_combout ;
wire \Selector0~13_combout ;
wire \Selector0~20_combout ;
wire \Selector0~14_combout ;
wire \Add1~1 ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~7 ;
wire \Add1~9 ;
wire \Add1~11 ;
wire \Add1~13 ;
wire \Add1~15 ;
wire \Add1~17 ;
wire \Add1~19 ;
wire \Add1~21 ;
wire \Add1~23 ;
wire \Add1~25 ;
wire \Add1~27 ;
wire \Add1~29 ;
wire \Add1~31 ;
wire \Add1~33 ;
wire \Add1~35 ;
wire \Add1~37 ;
wire \Add1~39 ;
wire \Add1~41 ;
wire \Add1~43 ;
wire \Add1~45 ;
wire \Add1~47 ;
wire \Add1~49 ;
wire \Add1~51 ;
wire \Add1~53 ;
wire \Add1~55 ;
wire \Add1~57 ;
wire \Add1~59 ;
wire \Add1~61 ;
wire \Add1~62_combout ;
wire \Selector0~17_combout ;
wire \Selector0~28_combout ;
wire \Selector0~15_combout ;
wire \Selector0~16_combout ;
wire \ShiftLeft0~12_combout ;
wire \ShiftLeft0~11_combout ;
wire \ShiftLeft0~13_combout ;
wire \ShiftLeft0~8_combout ;
wire \ShiftLeft0~9_combout ;
wire \Selector0~36_combout ;
wire \Selector1~9_combout ;
wire \Selector16~0_combout ;
wire \Selector0~23_combout ;
wire \Selector1~10_combout ;
wire \ShiftLeft0~15_combout ;
wire \ShiftLeft0~16_combout ;
wire \ShiftLeft0~17_combout ;
wire \Selector0~25_combout ;
wire \Selector0~26_combout ;
wire \Selector0~21_combout ;
wire \Selector0~29_combout ;
wire \Selector0~31_combout ;
wire \Add0~1 ;
wire \Add0~3 ;
wire \Add0~5 ;
wire \Add0~7 ;
wire \Add0~9 ;
wire \Add0~11 ;
wire \Add0~13 ;
wire \Add0~15 ;
wire \Add0~17 ;
wire \Add0~19 ;
wire \Add0~21 ;
wire \Add0~23 ;
wire \Add0~25 ;
wire \Add0~27 ;
wire \Add0~29 ;
wire \Add0~31 ;
wire \Add0~33 ;
wire \Add0~35 ;
wire \Add0~37 ;
wire \Add0~39 ;
wire \Add0~41 ;
wire \Add0~43 ;
wire \Add0~45 ;
wire \Add0~47 ;
wire \Add0~49 ;
wire \Add0~51 ;
wire \Add0~53 ;
wire \Add0~55 ;
wire \Add0~57 ;
wire \Add0~59 ;
wire \Add0~61 ;
wire \Add0~62_combout ;
wire \ShiftLeft0~22_combout ;
wire \ShiftLeft0~21_combout ;
wire \ShiftLeft0~18_combout ;
wire \ShiftLeft0~19_combout ;
wire \ShiftLeft0~20_combout ;
wire \ShiftLeft0~101_combout ;
wire \Selector1~8_combout ;
wire \Selector1~11_combout ;
wire \Selector0~30_combout ;
wire \Selector0~32_combout ;
wire \ShiftRight0~52_combout ;
wire \ShiftLeft0~43_combout ;
wire \ShiftLeft0~44_combout ;
wire \ShiftLeft0~45_combout ;
wire \Selector11~10_combout ;
wire \ShiftLeft0~40_combout ;
wire \ShiftLeft0~41_combout ;
wire \ShiftLeft0~42_combout ;
wire \ShiftLeft0~102_combout ;
wire \ShiftLeft0~48_combout ;
wire \Selector0~27_combout ;
wire \Selector3~1_combout ;
wire \Add0~56_combout ;
wire \Add1~56_combout ;
wire \Selector3~0_combout ;
wire \Selector3~2_combout ;
wire \ShiftRight0~124_combout ;
wire \Selector3~3_combout ;
wire \Selector0~18_combout ;
wire \Selector3~4_combout ;
wire \Selector3~5_combout ;
wire \Selector2~0_combout ;
wire \ShiftLeft0~29_combout ;
wire \ShiftLeft0~37_combout ;
wire \ShiftLeft0~33_combout ;
wire \ShiftLeft0~34_combout ;
wire \ShiftLeft0~35_combout ;
wire \ShiftLeft0~38_combout ;
wire \Selector3~6_combout ;
wire \ShiftRight0~51_combout ;
wire \ShiftLeft0~30_combout ;
wire \ShiftLeft0~31_combout ;
wire \Selector3~7_combout ;
wire \Selector3~8_combout ;
wire \Selector3~9_combout ;
wire \Selector7~14_combout ;
wire \Selector7~15_combout ;
wire \Selector7~16_combout ;
wire \Selector4~0_combout ;
wire \Selector7~8_combout ;
wire \Selector7~10_combout ;
wire \Selector7~18_combout ;
wire \ShiftLeft0~46_combout ;
wire \ShiftLeft0~47_combout ;
wire \ShiftLeft0~49_combout ;
wire \Selector7~11_combout ;
wire \ShiftLeft0~39_combout ;
wire \ShiftLeft0~50_combout ;
wire \ShiftLeft0~51_combout ;
wire \Selector7~12_combout ;
wire \Add1~48_combout ;
wire \Add0~48_combout ;
wire \Selector7~9_combout ;
wire \Selector7~13_combout ;
wire \Selector0~22_combout ;
wire \Selector8~2_combout ;
wire \Selector11~2_combout ;
wire \Selector11~4_combout ;
wire \Selector11~5_combout ;
wire \Selector11~6_combout ;
wire \Add1~40_combout ;
wire \Add0~40_combout ;
wire \Selector11~3_combout ;
wire \Selector11~7_combout ;
wire \Selector7~19_combout ;
wire \ShiftRight0~53_combout ;
wire \Selector15~0_combout ;
wire \Selector15~1_combout ;
wire \Selector15~3_combout ;
wire \Selector15~4_combout ;
wire \Selector15~5_combout ;
wire \Add0~32_combout ;
wire \Add1~32_combout ;
wire \Selector15~2_combout ;
wire \Selector15~6_combout ;
wire \Selector15~7_combout ;
wire \Selector28~1_combout ;
wire \Add1~6_combout ;
wire \Add0~6_combout ;
wire \Selector28~0_combout ;
wire \Selector28~2_combout ;
wire \Selector16~1_combout ;
wire \Selector28~3_combout ;
wire \Selector28~7_combout ;
wire \Selector28~4_combout ;
wire \ShiftRight0~55_combout ;
wire \ShiftRight0~62_combout ;
wire \ShiftRight0~60_combout ;
wire \ShiftRight0~61_combout ;
wire \ShiftRight0~63_combout ;
wire \ShiftRight0~64_combout ;
wire \ShiftRight0~59_combout ;
wire \ShiftRight0~57_combout ;
wire \ShiftRight0~58_combout ;
wire \Selector28~5_combout ;
wire \Selector28~6_combout ;
wire \Selector28~8_combout ;
wire \ShiftRight0~66_combout ;
wire \ShiftRight0~67_combout ;
wire \ShiftRight0~68_combout ;
wire \ShiftRight0~125_combout ;
wire \ShiftRight0~72_combout ;
wire \ShiftRight0~73_combout ;
wire \ShiftRight0~69_combout ;
wire \ShiftRight0~70_combout ;
wire \ShiftRight0~71_combout ;
wire \Selector20~0_combout ;
wire \ShiftRight0~74_combout ;
wire \ShiftLeft0~52_combout ;
wire \ShiftLeft0~53_combout ;
wire \Selector29~0_combout ;
wire \Selector29~2_combout ;
wire \Add1~4_combout ;
wire \Add0~4_combout ;
wire \Selector29~1_combout ;
wire \Selector29~3_combout ;
wire \ShiftRight0~80_combout ;
wire \ShiftRight0~77_combout ;
wire \ShiftRight0~78_combout ;
wire \ShiftRight0~81_combout ;
wire \ShiftRight0~41_combout ;
wire \ShiftRight0~75_combout ;
wire \ShiftRight0~76_combout ;
wire \Selector29~4_combout ;
wire \Selector29~5_combout ;
wire \Selector29~6_combout ;
wire \ShiftRight0~83_combout ;
wire \ShiftRight0~82_combout ;
wire \ShiftRight0~84_combout ;
wire \ShiftRight0~88_combout ;
wire \ShiftRight0~86_combout ;
wire \ShiftRight0~87_combout ;
wire \ShiftRight0~89_combout ;
wire \Selector21~0_combout ;
wire \ShiftLeft0~55_combout ;
wire \ShiftLeft0~54_combout ;
wire \ShiftLeft0~56_combout ;
wire \ShiftLeft0~61_combout ;
wire \ShiftLeft0~58_combout ;
wire \ShiftLeft0~59_combout ;
wire \ShiftLeft0~60_combout ;
wire \Selector10~0_combout ;
wire \Add1~42_combout ;
wire \Add0~42_combout ;
wire \Selector10~2_combout ;
wire \Selector10~3_combout ;
wire \Selector10~4_combout ;
wire \Selector10~5_combout ;
wire \ShiftRight0~97_combout ;
wire \ShiftRight0~98_combout ;
wire \ShiftRight0~94_combout ;
wire \ShiftRight0~95_combout ;
wire \ShiftRight0~96_combout ;
wire \ShiftRight0~99_combout ;
wire \ShiftLeft0~63_combout ;
wire \ShiftLeft0~66_combout ;
wire \ShiftLeft0~65_combout ;
wire \ShiftLeft0~67_combout ;
wire \ShiftLeft0~62_combout ;
wire \ShiftLeft0~103_combout ;
wire \Selector2~7_combout ;
wire \Selector2~8_combout ;
wire \Add1~58_combout ;
wire \ShiftLeft0~68_combout ;
wire \ShiftLeft0~69_combout ;
wire \ShiftLeft0~70_combout ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \Selector2~5_combout ;
wire \Selector2~3_combout ;
wire \Add0~58_combout ;
wire \Selector2~4_combout ;
wire \Selector2~6_combout ;
wire \Selector1~16_combout ;
wire \Add0~60_combout ;
wire \Selector1~17_combout ;
wire \Selector1~18_combout ;
wire \ShiftLeft0~71_combout ;
wire \ShiftLeft0~72_combout ;
wire \ShiftLeft0~73_combout ;
wire \ShiftLeft0~74_combout ;
wire \ShiftLeft0~75_combout ;
wire \ShiftLeft0~76_combout ;
wire \ShiftLeft0~77_combout ;
wire \ShiftLeft0~79_combout ;
wire \ShiftLeft0~78_combout ;
wire \Selector9~0_combout ;
wire \Selector1~12_combout ;
wire \Selector1~22_combout ;
wire \Add1~60_combout ;
wire \Selector1~20_combout ;
wire \Selector1~19_combout ;
wire \Selector1~21_combout ;
wire \Selector1~23_combout ;
wire \ShiftLeft0~32_combout ;
wire \Selector1~13_combout ;
wire \ShiftLeft0~80_combout ;
wire \ShiftLeft0~81_combout ;
wire \Selector1~14_combout ;
wire \Selector1~15_combout ;
wire \Selector0~7_combout ;
wire \Selector4~7_combout ;
wire \Selector4~8_combout ;
wire \Selector4~9_combout ;
wire \ShiftLeft0~24_combout ;
wire \ShiftLeft0~26_combout ;
wire \ShiftLeft0~89_combout ;
wire \ShiftLeft0~90_combout ;
wire \Selector4~4_combout ;
wire \Selector4~5_combout ;
wire \Add1~54_combout ;
wire \Add0~54_combout ;
wire \Selector4~2_combout ;
wire \Selector4~3_combout ;
wire \Selector4~6_combout ;
wire \Selector5~2_combout ;
wire \Selector5~3_combout ;
wire \Selector5~4_combout ;
wire \ShiftLeft0~92_combout ;
wire \ShiftLeft0~93_combout ;
wire \ShiftLeft0~86_combout ;
wire \ShiftLeft0~85_combout ;
wire \ShiftLeft0~87_combout ;
wire \ShiftLeft0~82_combout ;
wire \ShiftLeft0~83_combout ;
wire \ShiftLeft0~84_combout ;
wire \ShiftLeft0~91_combout ;
wire \Selector5~5_combout ;
wire \Selector5~6_combout ;
wire \Add1~52_combout ;
wire \Add0~52_combout ;
wire \Selector5~0_combout ;
wire \Selector5~1_combout ;
wire \ShiftLeft0~23_combout ;
wire \Selector12~0_combout ;
wire \Selector12~1_combout ;
wire \ShiftLeft0~10_combout ;
wire \ShiftLeft0~28_combout ;
wire \ShiftLeft0~27_combout ;
wire \ShiftLeft0~88_combout ;
wire \Add1~38_combout ;
wire \Add0~38_combout ;
wire \Selector12~2_combout ;
wire \Selector12~6_combout ;
wire \Selector12~7_combout ;
wire \Selector24~6_combout ;
wire \Selector24~7_combout ;
wire \Selector24~8_combout ;
wire \Add0~14_combout ;
wire \Add1~14_combout ;
wire \Selector24~2_combout ;
wire \Selector24~1_combout ;
wire \ShiftRight0~100_combout ;
wire \Selector24~3_combout ;
wire \ShiftRight0~65_combout ;
wire \ShiftRight0~102_combout ;
wire \ShiftRight0~103_combout ;
wire \Selector24~4_combout ;
wire \Selector24~5_combout ;
wire \Selector13~0_combout ;
wire \Selector13~1_combout ;
wire \Add1~36_combout ;
wire \Add0~36_combout ;
wire \Selector13~2_combout ;
wire \Selector13~6_combout ;
wire \Selector13~7_combout ;
wire \Selector25~5_combout ;
wire \Selector25~6_combout ;
wire \Selector25~7_combout ;
wire \Selector25~0_combout ;
wire \Selector0~10_combout ;
wire \Add0~12_combout ;
wire \Add1~12_combout ;
wire \Selector25~1_combout ;
wire \ShiftRight0~105_combout ;
wire \Selector25~2_combout ;
wire \ShiftRight0~107_combout ;
wire \ShiftRight0~108_combout ;
wire \Selector25~3_combout ;
wire \Selector25~4_combout ;
wire \Selector1~25_combout ;
wire \ShiftLeft0~94_combout ;
wire \Selector14~0_combout ;
wire \Selector14~3_combout ;
wire \Selector14~4_combout ;
wire \Selector14~5_combout ;
wire \Add1~34_combout ;
wire \Add0~34_combout ;
wire \Selector14~2_combout ;
wire \ShiftLeft0~64_combout ;
wire \ShiftLeft0~95_combout ;
wire \ShiftRight0~92_combout ;
wire \ShiftRight0~91_combout ;
wire \ShiftRight0~93_combout ;
wire \ShiftRight0~109_combout ;
wire \ShiftRight0~110_combout ;
wire \ShiftRight0~111_combout ;
wire \Selector22~1_combout ;
wire \ShiftRight0~112_combout ;
wire \Selector27~5_combout ;
wire \Selector27~6_combout ;
wire \Selector27~7_combout ;
wire \Add0~8_combout ;
wire \Add1~8_combout ;
wire \Selector27~0_combout ;
wire \Selector27~1_combout ;
wire \Selector27~3_combout ;
wire \Selector27~4_combout ;
wire \Selector8~1_combout ;
wire \ShiftLeft0~96_combout ;
wire \Selector16~3_combout ;
wire \Selector16~4_combout ;
wire \Selector16~5_combout ;
wire \Add1~30_combout ;
wire \Add0~30_combout ;
wire \Selector16~2_combout ;
wire \Selector16~6_combout ;
wire \Selector16~9_combout ;
wire \Selector16~8_combout ;
wire \Selector0~35_combout ;
wire \Selector16~7_combout ;
wire \Selector16~10_combout ;
wire \Selector18~0_combout ;
wire \Selector18~1_combout ;
wire \Add0~26_combout ;
wire \Selector18~2_combout ;
wire \Selector18~6_combout ;
wire \ShiftRight0~115_combout ;
wire \ShiftRight0~114_combout ;
wire \ShiftRight0~116_combout ;
wire \Selector18~7_combout ;
wire \ShiftLeft0~97_combout ;
wire \ShiftLeft0~98_combout ;
wire \Selector17~0_combout ;
wire \Selector17~1_combout ;
wire \ShiftRight0~106_combout ;
wire \Add1~28_combout ;
wire \Add0~28_combout ;
wire \Selector17~2_combout ;
wire \Selector17~6_combout ;
wire \Selector17~7_combout ;
wire \Selector6~2_combout ;
wire \Selector6~5_combout ;
wire \Add1~50_combout ;
wire \Add0~50_combout ;
wire \Selector6~3_combout ;
wire \Selector6~4_combout ;
wire \Selector6~6_combout ;
wire \Selector6~0_combout ;
wire \ShiftLeft0~99_combout ;
wire \ShiftLeft0~100_combout ;
wire \Selector6~1_combout ;
wire \Add0~10_combout ;
wire \Add1~10_combout ;
wire \Selector26~0_combout ;
wire \Selector26~1_combout ;
wire \Selector26~2_combout ;
wire \Selector26~3_combout ;
wire \Selector26~4_combout ;
wire \ShiftRight0~119_combout ;
wire \ShiftRight0~120_combout ;
wire \ShiftRight0~117_combout ;
wire \ShiftRight0~118_combout ;
wire \Selector26~5_combout ;
wire \Selector26~6_combout ;
wire \Selector19~0_combout ;
wire \Selector19~1_combout ;
wire \ShiftRight0~34_combout ;
wire \ShiftRight0~113_combout ;
wire \Selector19~4_combout ;
wire \Selector19~5_combout ;
wire \Selector19~6_combout ;
wire \Add1~24_combout ;
wire \Add0~24_combout ;
wire \Selector19~2_combout ;
wire \Selector19~3_combout ;
wire \Selector19~7_combout ;
wire \Selector20~1_combout ;
wire \Add0~22_combout ;
wire \Add1~22_combout ;
wire \Selector20~3_combout ;
wire \Selector20~4_combout ;
wire \Selector20~5_combout ;
wire \Selector20~6_combout ;
wire \Selector21~3_combout ;
wire \Selector21~4_combout ;
wire \Selector21~5_combout ;
wire \Add1~20_combout ;
wire \Add0~20_combout ;
wire \Selector21~2_combout ;
wire \Selector8~5_combout ;
wire \Selector8~6_combout ;
wire \Selector8~7_combout ;
wire \Add1~46_combout ;
wire \Add0~46_combout ;
wire \Selector8~4_combout ;
wire \Selector9~3_combout ;
wire \Selector9~4_combout ;
wire \Selector9~5_combout ;
wire \Add1~44_combout ;
wire \Add0~44_combout ;
wire \Selector9~2_combout ;
wire \Selector1~26_combout ;
wire \Selector22~2_combout ;
wire \Selector22~5_combout ;
wire \Selector22~6_combout ;
wire \Selector22~7_combout ;
wire \Add1~18_combout ;
wire \Add0~18_combout ;
wire \Selector22~3_combout ;
wire \Selector22~4_combout ;
wire \Selector30~2_combout ;
wire \Selector22~8_combout ;
wire \Selector30~8_combout ;
wire \Selector30~3_combout ;
wire \Selector30~4_combout ;
wire \Add1~2_combout ;
wire \Selector30~5_combout ;
wire \Selector30~6_combout ;
wire \Selector30~7_combout ;
wire \Selector30~15_combout ;
wire \Selector30~9_combout ;
wire \Selector30~11_combout ;
wire \Selector30~12_combout ;
wire \Selector30~10_combout ;
wire \Selector30~13_combout ;
wire \ShiftRight0~121_combout ;
wire \Selector23~6_combout ;
wire \Selector23~7_combout ;
wire \Selector23~8_combout ;
wire \Add0~16_combout ;
wire \Add1~16_combout ;
wire \Selector23~5_combout ;
wire \Selector23~9_combout ;
wire \Equal0~2_combout ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~3_combout ;
wire \Equal0~10_combout ;
wire \Equal0~5_combout ;
wire \Equal0~7_combout ;
wire \Equal0~4_combout ;
wire \Equal0~6_combout ;
wire \Equal0~8_combout ;
wire \Equal0~9_combout ;


// Location: LCCOMB_X56_Y37_N26
cycloneive_lcell_comb \Add1~26 (
// Equation(s):
// \Add1~26_combout  = (\portB~39_combout  & ((Mux18 & (!\Add1~25 )) # (!Mux18 & ((\Add1~25 ) # (GND))))) # (!\portB~39_combout  & ((Mux18 & (\Add1~25  & VCC)) # (!Mux18 & (!\Add1~25 ))))
// \Add1~27  = CARRY((\portB~39_combout  & ((!\Add1~25 ) # (!Mux18))) # (!\portB~39_combout  & (!Mux18 & !\Add1~25 )))

	.dataa(portB18),
	.datab(Mux18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~25 ),
	.combout(\Add1~26_combout ),
	.cout(\Add1~27 ));
// synopsys translate_off
defparam \Add1~26 .lut_mask = 16'h692B;
defparam \Add1~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N2
cycloneive_lcell_comb \Add0~2 (
// Equation(s):
// \Add0~2_combout  = (\portB~63_combout  & ((Mux302 & (\Add0~1  & VCC)) # (!Mux302 & (!\Add0~1 )))) # (!\portB~63_combout  & ((Mux302 & (!\Add0~1 )) # (!Mux302 & ((\Add0~1 ) # (GND)))))
// \Add0~3  = CARRY((\portB~63_combout  & (!Mux302 & !\Add0~1 )) # (!\portB~63_combout  & ((!\Add0~1 ) # (!Mux302))))

	.dataa(portB30),
	.datab(Mux302),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
// synopsys translate_off
defparam \Add0~2 .lut_mask = 16'h9617;
defparam \Add0~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N18
cycloneive_lcell_comb \ShiftRight0~15 (
// Equation(s):
// \ShiftRight0~15_combout  = (Mux5) # ((Mux4) # ((Mux6) # (Mux72)))

	.dataa(Mux5),
	.datab(Mux4),
	.datac(Mux6),
	.datad(Mux72),
	.cin(gnd),
	.combout(\ShiftRight0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~15 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N2
cycloneive_lcell_comb \ShiftRight0~21 (
// Equation(s):
// \ShiftRight0~21_combout  = (Mux26) # ((Mux242) # (Mux252))

	.dataa(Mux26),
	.datab(Mux242),
	.datac(gnd),
	.datad(Mux252),
	.cin(gnd),
	.combout(\ShiftRight0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~21 .lut_mask = 16'hFFEE;
defparam \ShiftRight0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N22
cycloneive_lcell_comb \Selector0~19 (
// Equation(s):
// \Selector0~19_combout  = (\Selector0~17_combout ) # ((\Selector0~18_combout  & Mux0))

	.dataa(\Selector0~18_combout ),
	.datab(gnd),
	.datac(\Selector0~17_combout ),
	.datad(Mux0),
	.cin(gnd),
	.combout(\Selector0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~19 .lut_mask = 16'hFAF0;
defparam \Selector0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N6
cycloneive_lcell_comb \ShiftLeft0~14 (
// Equation(s):
// \ShiftLeft0~14_combout  = (Mux312 & ((\portB~9_combout ))) # (!Mux312 & (\portB~7_combout ))

	.dataa(gnd),
	.datab(portB2),
	.datac(Mux312),
	.datad(portB3),
	.cin(gnd),
	.combout(\ShiftLeft0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~14 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N26
cycloneive_lcell_comb \Selector0~24 (
// Equation(s):
// \Selector0~24_combout  = (\Selector1~25_combout  & (((\Selector1~10_combout ) # (\ShiftLeft0~14_combout )))) # (!\Selector1~25_combout  & (\portB~3_combout  & (!\Selector1~10_combout )))

	.dataa(\Selector1~25_combout ),
	.datab(portB),
	.datac(\Selector1~10_combout ),
	.datad(\ShiftLeft0~14_combout ),
	.cin(gnd),
	.combout(\Selector0~24_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~24 .lut_mask = 16'hAEA4;
defparam \Selector0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N30
cycloneive_lcell_comb \ShiftLeft0~25 (
// Equation(s):
// \ShiftLeft0~25_combout  = (\portB~47_combout  & ((\ShiftRight0~122_combout ) # ((\portB~43_combout  & \ShiftRight0~123_combout )))) # (!\portB~47_combout  & (((\portB~43_combout  & \ShiftRight0~123_combout ))))

	.dataa(portB22),
	.datab(\ShiftRight0~122_combout ),
	.datac(portB20),
	.datad(\ShiftRight0~123_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~25 .lut_mask = 16'hF888;
defparam \ShiftLeft0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N14
cycloneive_lcell_comb \ShiftLeft0~36 (
// Equation(s):
// \ShiftLeft0~36_combout  = (Mux312 & ((Mux302 & ((\portB~39_combout ))) # (!Mux302 & (\portB~35_combout ))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB16),
	.datad(portB18),
	.cin(gnd),
	.combout(\ShiftLeft0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~36 .lut_mask = 16'hA820;
defparam \ShiftLeft0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N6
cycloneive_lcell_comb \Selector0~34 (
// Equation(s):
// \Selector0~34_combout  = (!cuifALUOP_2 & (!cuifALUOP_1 & (!cuifALUOP_0 & !cuifALUOP_3)))

	.dataa(cuifALUOP_2),
	.datab(cuifALUOP_1),
	.datac(cuifALUOP_0),
	.datad(cuifALUOP_3),
	.cin(gnd),
	.combout(\Selector0~34_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~34 .lut_mask = 16'h0001;
defparam \Selector0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N12
cycloneive_lcell_comb \ShiftRight0~56 (
// Equation(s):
// \ShiftRight0~56_combout  = (Mux312 & (\portB~49_combout  & !Mux302))

	.dataa(Mux312),
	.datab(portB23),
	.datac(gnd),
	.datad(Mux302),
	.cin(gnd),
	.combout(\ShiftRight0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~56 .lut_mask = 16'h0088;
defparam \ShiftRight0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N14
cycloneive_lcell_comb \ShiftRight0~79 (
// Equation(s):
// \ShiftRight0~79_combout  = (!Mux302 & ((Mux312 & (\portB~43_combout )) # (!Mux312 & ((\portB~45_combout )))))

	.dataa(portB20),
	.datab(portB21),
	.datac(Mux302),
	.datad(Mux312),
	.cin(gnd),
	.combout(\ShiftRight0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~79 .lut_mask = 16'h0A0C;
defparam \ShiftRight0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N14
cycloneive_lcell_comb \Selector12~3 (
// Equation(s):
// \Selector12~3_combout  = (\portB~27_combout  & ((\Selector0~17_combout ) # ((Mux12 & \Selector0~18_combout ))))

	.dataa(portB12),
	.datab(\Selector0~17_combout ),
	.datac(Mux12),
	.datad(\Selector0~18_combout ),
	.cin(gnd),
	.combout(\Selector12~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~3 .lut_mask = 16'hA888;
defparam \Selector12~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N8
cycloneive_lcell_comb \Selector12~4 (
// Equation(s):
// \Selector12~4_combout  = (\Selector12~3_combout ) # ((\Selector0~27_combout  & (!Mux12 & !\portB~27_combout )))

	.dataa(\Selector0~27_combout ),
	.datab(\Selector12~3_combout ),
	.datac(Mux12),
	.datad(portB12),
	.cin(gnd),
	.combout(\Selector12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~4 .lut_mask = 16'hCCCE;
defparam \Selector12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N26
cycloneive_lcell_comb \Selector12~5 (
// Equation(s):
// \Selector12~5_combout  = (\Selector12~4_combout ) # ((\Selector0~15_combout  & (\portB~27_combout  $ (Mux12))))

	.dataa(portB12),
	.datab(\Selector12~4_combout ),
	.datac(Mux12),
	.datad(\Selector0~15_combout ),
	.cin(gnd),
	.combout(\Selector12~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~5 .lut_mask = 16'hDECC;
defparam \Selector12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N30
cycloneive_lcell_comb \ShiftRight0~101 (
// Equation(s):
// \ShiftRight0~101_combout  = (\ShiftRight0~62_combout ) # (\ShiftRight0~63_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftRight0~62_combout ),
	.datad(\ShiftRight0~63_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~101_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~101 .lut_mask = 16'hFFF0;
defparam \ShiftRight0~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N6
cycloneive_lcell_comb \Selector13~3 (
// Equation(s):
// \Selector13~3_combout  = (\portB~29_combout  & ((\Selector0~17_combout ) # ((\Selector0~18_combout  & Mux13))))

	.dataa(\Selector0~18_combout ),
	.datab(Mux13),
	.datac(\Selector0~17_combout ),
	.datad(portB13),
	.cin(gnd),
	.combout(\Selector13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~3 .lut_mask = 16'hF800;
defparam \Selector13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N8
cycloneive_lcell_comb \Selector13~4 (
// Equation(s):
// \Selector13~4_combout  = (\Selector13~3_combout ) # ((!\portB~29_combout  & (!Mux13 & \Selector0~27_combout )))

	.dataa(\Selector13~3_combout ),
	.datab(portB13),
	.datac(Mux13),
	.datad(\Selector0~27_combout ),
	.cin(gnd),
	.combout(\Selector13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~4 .lut_mask = 16'hABAA;
defparam \Selector13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N26
cycloneive_lcell_comb \Selector13~5 (
// Equation(s):
// \Selector13~5_combout  = (\Selector13~4_combout ) # ((\Selector0~15_combout  & (Mux13 $ (\portB~29_combout ))))

	.dataa(Mux13),
	.datab(portB13),
	.datac(\Selector13~4_combout ),
	.datad(\Selector0~15_combout ),
	.cin(gnd),
	.combout(\Selector13~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~5 .lut_mask = 16'hF6F0;
defparam \Selector13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N30
cycloneive_lcell_comb \ShiftRight0~104 (
// Equation(s):
// \ShiftRight0~104_combout  = (\ShiftRight0~80_combout ) # (\ShiftRight0~79_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftRight0~80_combout ),
	.datad(\ShiftRight0~79_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~104_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~104 .lut_mask = 16'hFFF0;
defparam \ShiftRight0~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N22
cycloneive_lcell_comb \Selector27~2 (
// Equation(s):
// \Selector27~2_combout  = (\Selector7~18_combout  & ((\Selector7~10_combout ) # ((\ShiftRight0~113_combout )))) # (!\Selector7~18_combout  & (!\Selector7~10_combout  & ((\ShiftRight0~42_combout ))))

	.dataa(\Selector7~18_combout ),
	.datab(\Selector7~10_combout ),
	.datac(\ShiftRight0~113_combout ),
	.datad(\ShiftRight0~42_combout ),
	.cin(gnd),
	.combout(\Selector27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~2 .lut_mask = 16'hB9A8;
defparam \Selector27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N28
cycloneive_lcell_comb \Selector18~3 (
// Equation(s):
// \Selector18~3_combout  = (\portB~39_combout  & ((\Selector0~17_combout ) # ((\Selector0~18_combout  & Mux18))))

	.dataa(\Selector0~18_combout ),
	.datab(portB18),
	.datac(Mux18),
	.datad(\Selector0~17_combout ),
	.cin(gnd),
	.combout(\Selector18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~3 .lut_mask = 16'hCC80;
defparam \Selector18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N26
cycloneive_lcell_comb \Selector18~4 (
// Equation(s):
// \Selector18~4_combout  = (\Selector18~3_combout ) # ((\Selector0~27_combout  & (!\portB~39_combout  & !Mux18)))

	.dataa(\Selector0~27_combout ),
	.datab(portB18),
	.datac(Mux18),
	.datad(\Selector18~3_combout ),
	.cin(gnd),
	.combout(\Selector18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~4 .lut_mask = 16'hFF02;
defparam \Selector18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N12
cycloneive_lcell_comb \Selector18~5 (
// Equation(s):
// \Selector18~5_combout  = (\Selector18~4_combout ) # ((\Selector0~15_combout  & (\portB~39_combout  $ (Mux18))))

	.dataa(portB18),
	.datab(Mux18),
	.datac(\Selector18~4_combout ),
	.datad(\Selector0~15_combout ),
	.cin(gnd),
	.combout(\Selector18~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~5 .lut_mask = 16'hF6F0;
defparam \Selector18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N0
cycloneive_lcell_comb \Selector17~3 (
// Equation(s):
// \Selector17~3_combout  = (\portB~37_combout  & ((\Selector0~17_combout ) # ((\Selector0~18_combout  & Mux17))))

	.dataa(\Selector0~18_combout ),
	.datab(\Selector0~17_combout ),
	.datac(Mux17),
	.datad(portB17),
	.cin(gnd),
	.combout(\Selector17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~3 .lut_mask = 16'hEC00;
defparam \Selector17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N2
cycloneive_lcell_comb \Selector17~4 (
// Equation(s):
// \Selector17~4_combout  = (\Selector17~3_combout ) # ((\Selector0~27_combout  & (!\portB~37_combout  & !Mux17)))

	.dataa(\Selector0~27_combout ),
	.datab(portB17),
	.datac(Mux17),
	.datad(\Selector17~3_combout ),
	.cin(gnd),
	.combout(\Selector17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~4 .lut_mask = 16'hFF02;
defparam \Selector17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N4
cycloneive_lcell_comb \Selector17~5 (
// Equation(s):
// \Selector17~5_combout  = (\Selector17~4_combout ) # ((\Selector0~15_combout  & (Mux17 $ (\portB~37_combout ))))

	.dataa(\Selector0~15_combout ),
	.datab(\Selector17~4_combout ),
	.datac(Mux17),
	.datad(portB17),
	.cin(gnd),
	.combout(\Selector17~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~5 .lut_mask = 16'hCEEC;
defparam \Selector17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N20
cycloneive_lcell_comb \Selector31~10 (
// Equation(s):
// Selector31 = (\Selector31~7_combout ) # ((\Selector31~9_combout ) # ((\Selector0~4_combout  & \LessThan1~62_combout )))

	.dataa(\Selector0~4_combout ),
	.datab(\Selector31~7_combout ),
	.datac(\Selector31~9_combout ),
	.datad(\LessThan1~62_combout ),
	.cin(gnd),
	.combout(Selector31),
	.cout());
// synopsys translate_off
defparam \Selector31~10 .lut_mask = 16'hFEFC;
defparam \Selector31~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N12
cycloneive_lcell_comb \ShiftRight0~50 (
// Equation(s):
// ShiftRight0 = (Mux272 & (((\ShiftRight0~36_combout )))) # (!Mux272 & ((\ShiftRight0~43_combout ) # ((\ShiftRight0~49_combout ))))

	.dataa(Mux272),
	.datab(\ShiftRight0~43_combout ),
	.datac(\ShiftRight0~49_combout ),
	.datad(\ShiftRight0~36_combout ),
	.cin(gnd),
	.combout(ShiftRight0),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~50 .lut_mask = 16'hFE54;
defparam \ShiftRight0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N22
cycloneive_lcell_comb \Selector24~0 (
// Equation(s):
// Selector24 = (\Selector0~13_combout  & !\ShiftRight0~22_combout )

	.dataa(\Selector0~13_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ShiftRight0~22_combout ),
	.cin(gnd),
	.combout(Selector24),
	.cout());
// synopsys translate_off
defparam \Selector24~0 .lut_mask = 16'h00AA;
defparam \Selector24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N22
cycloneive_lcell_comb \Selector8~0 (
// Equation(s):
// Selector8 = (!Mux272 & (\Selector0~20_combout  & !\ShiftRight0~22_combout ))

	.dataa(gnd),
	.datab(Mux272),
	.datac(\Selector0~20_combout ),
	.datad(\ShiftRight0~22_combout ),
	.cin(gnd),
	.combout(Selector8),
	.cout());
// synopsys translate_off
defparam \Selector8~0 .lut_mask = 16'h0030;
defparam \Selector8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N6
cycloneive_lcell_comb \Selector0~33 (
// Equation(s):
// Selector0 = (\Selector0~29_combout ) # ((\Selector0~32_combout ) # ((\Selector0~14_combout  & \Add1~62_combout )))

	.dataa(\Selector0~14_combout ),
	.datab(\Add1~62_combout ),
	.datac(\Selector0~29_combout ),
	.datad(\Selector0~32_combout ),
	.cin(gnd),
	.combout(Selector0),
	.cout());
// synopsys translate_off
defparam \Selector0~33 .lut_mask = 16'hFFF8;
defparam \Selector0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N6
cycloneive_lcell_comb \Selector3~10 (
// Equation(s):
// Selector3 = (\Selector3~2_combout ) # ((\Selector3~9_combout ) # ((\Selector1~11_combout  & \ShiftLeft0~48_combout )))

	.dataa(\Selector1~11_combout ),
	.datab(\ShiftLeft0~48_combout ),
	.datac(\Selector3~2_combout ),
	.datad(\Selector3~9_combout ),
	.cin(gnd),
	.combout(Selector3),
	.cout());
// synopsys translate_off
defparam \Selector3~10 .lut_mask = 16'hFFF8;
defparam \Selector3~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N4
cycloneive_lcell_comb \Selector4~1 (
// Equation(s):
// Selector4 = (!Mux28 & (\Selector0~13_combout  & (!Mux272 & !\ShiftRight0~22_combout )))

	.dataa(Mux28),
	.datab(\Selector0~13_combout ),
	.datac(Mux272),
	.datad(\ShiftRight0~22_combout ),
	.cin(gnd),
	.combout(Selector4),
	.cout());
// synopsys translate_off
defparam \Selector4~1 .lut_mask = 16'h0004;
defparam \Selector4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N30
cycloneive_lcell_comb \Selector7~17 (
// Equation(s):
// Selector7 = (\Selector7~16_combout ) # ((\Selector7~13_combout ) # ((Selector4 & \ShiftRight0~30_combout )))

	.dataa(Selector4),
	.datab(\ShiftRight0~30_combout ),
	.datac(\Selector7~16_combout ),
	.datad(\Selector7~13_combout ),
	.cin(gnd),
	.combout(Selector7),
	.cout());
// synopsys translate_off
defparam \Selector7~17 .lut_mask = 16'hFFF8;
defparam \Selector7~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N10
cycloneive_lcell_comb \Selector11~8 (
// Equation(s):
// Selector11 = (\Selector11~2_combout ) # ((\Selector11~7_combout ) # ((\Selector0~23_combout  & \ShiftLeft0~38_combout )))

	.dataa(\Selector0~23_combout ),
	.datab(\Selector11~2_combout ),
	.datac(\ShiftLeft0~38_combout ),
	.datad(\Selector11~7_combout ),
	.cin(gnd),
	.combout(Selector11),
	.cout());
// synopsys translate_off
defparam \Selector11~8 .lut_mask = 16'hFFEC;
defparam \Selector11~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N4
cycloneive_lcell_comb \ShiftRight0~54 (
// Equation(s):
// ShiftRight01 = (\ShiftRight0~53_combout ) # ((Mux28 & (\ShiftRight0~26_combout  & !Mux292)))

	.dataa(Mux28),
	.datab(\ShiftRight0~26_combout ),
	.datac(Mux292),
	.datad(\ShiftRight0~53_combout ),
	.cin(gnd),
	.combout(ShiftRight01),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~54 .lut_mask = 16'hFF08;
defparam \ShiftRight0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N30
cycloneive_lcell_comb \Selector11~9 (
// Equation(s):
// Selector111 = (Selector11) # ((Selector8 & ShiftRight01))

	.dataa(gnd),
	.datab(Selector8),
	.datac(ShiftRight01),
	.datad(Selector11),
	.cin(gnd),
	.combout(Selector111),
	.cout());
// synopsys translate_off
defparam \Selector11~9 .lut_mask = 16'hFFC0;
defparam \Selector11~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N12
cycloneive_lcell_comb \Selector15~8 (
// Equation(s):
// Selector15 = (\Selector15~1_combout ) # ((\Selector15~7_combout ) # ((Selector8 & \ShiftRight0~36_combout )))

	.dataa(Selector8),
	.datab(\ShiftRight0~36_combout ),
	.datac(\Selector15~1_combout ),
	.datad(\Selector15~7_combout ),
	.cin(gnd),
	.combout(Selector15),
	.cout());
// synopsys translate_off
defparam \Selector15~8 .lut_mask = 16'hFFF8;
defparam \Selector15~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N10
cycloneive_lcell_comb \Selector22~0 (
// Equation(s):
// Selector22 = (cuifALUOP_0 & (Mux272 & \Selector1~8_combout ))

	.dataa(cuifALUOP_0),
	.datab(Mux272),
	.datac(gnd),
	.datad(\Selector1~8_combout ),
	.cin(gnd),
	.combout(Selector22),
	.cout());
// synopsys translate_off
defparam \Selector22~0 .lut_mask = 16'h8800;
defparam \Selector22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N4
cycloneive_lcell_comb \Selector28~9 (
// Equation(s):
// Selector28 = (\Selector28~2_combout ) # ((\Selector28~8_combout ) # ((Selector22 & \ShiftRight0~74_combout )))

	.dataa(\Selector28~2_combout ),
	.datab(Selector22),
	.datac(\Selector28~8_combout ),
	.datad(\ShiftRight0~74_combout ),
	.cin(gnd),
	.combout(Selector28),
	.cout());
// synopsys translate_off
defparam \Selector28~9 .lut_mask = 16'hFEFA;
defparam \Selector28~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N8
cycloneive_lcell_comb \Selector29~7 (
// Equation(s):
// Selector29 = (\Selector29~6_combout ) # ((\ShiftLeft0~53_combout  & (\ShiftRight0~124_combout  & \Selector16~1_combout )))

	.dataa(\ShiftLeft0~53_combout ),
	.datab(\Selector29~6_combout ),
	.datac(\ShiftRight0~124_combout ),
	.datad(\Selector16~1_combout ),
	.cin(gnd),
	.combout(Selector29),
	.cout());
// synopsys translate_off
defparam \Selector29~7 .lut_mask = 16'hECCC;
defparam \Selector29~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N14
cycloneive_lcell_comb \ShiftRight0~85 (
// Equation(s):
// ShiftRight02 = (Mux292 & (((!Mux302 & \ShiftRight0~25_combout )))) # (!Mux292 & (\ShiftRight0~84_combout ))

	.dataa(Mux292),
	.datab(\ShiftRight0~84_combout ),
	.datac(Mux302),
	.datad(\ShiftRight0~25_combout ),
	.cin(gnd),
	.combout(ShiftRight02),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~85 .lut_mask = 16'h4E44;
defparam \ShiftRight0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N30
cycloneive_lcell_comb \ShiftRight0~90 (
// Equation(s):
// ShiftRight03 = (Mux28 & ((ShiftRight02))) # (!Mux28 & (\Selector21~0_combout ))

	.dataa(gnd),
	.datab(Mux28),
	.datac(\Selector21~0_combout ),
	.datad(ShiftRight02),
	.cin(gnd),
	.combout(ShiftRight03),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~90 .lut_mask = 16'hFC30;
defparam \ShiftRight0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N26
cycloneive_lcell_comb \Selector29~8 (
// Equation(s):
// Selector291 = (Selector29) # ((Selector22 & ShiftRight03))

	.dataa(gnd),
	.datab(Selector22),
	.datac(Selector29),
	.datad(ShiftRight03),
	.cin(gnd),
	.combout(Selector291),
	.cout());
// synopsys translate_off
defparam \Selector29~8 .lut_mask = 16'hFCF0;
defparam \Selector29~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N18
cycloneive_lcell_comb \ShiftLeft0~57 (
// Equation(s):
// ShiftLeft0 = (\ShiftLeft0~56_combout ) # ((Mux292 & (!Mux302 & \ShiftLeft0~19_combout )))

	.dataa(Mux292),
	.datab(Mux302),
	.datac(\ShiftLeft0~56_combout ),
	.datad(\ShiftLeft0~19_combout ),
	.cin(gnd),
	.combout(ShiftLeft0),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~57 .lut_mask = 16'hF2F0;
defparam \ShiftLeft0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N26
cycloneive_lcell_comb \Selector10~1 (
// Equation(s):
// Selector10 = (\Selector8~2_combout  & ((ShiftLeft0) # ((\Selector0~22_combout  & \Selector10~0_combout )))) # (!\Selector8~2_combout  & (\Selector0~22_combout  & (\Selector10~0_combout )))

	.dataa(\Selector8~2_combout ),
	.datab(\Selector0~22_combout ),
	.datac(\Selector10~0_combout ),
	.datad(ShiftLeft0),
	.cin(gnd),
	.combout(Selector10),
	.cout());
// synopsys translate_off
defparam \Selector10~1 .lut_mask = 16'hEAC0;
defparam \Selector10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N28
cycloneive_lcell_comb \Selector10~6 (
// Equation(s):
// Selector101 = (\Selector10~2_combout ) # ((\Selector10~5_combout ) # ((Mux10 & \Selector0~17_combout )))

	.dataa(Mux10),
	.datab(\Selector0~17_combout ),
	.datac(\Selector10~2_combout ),
	.datad(\Selector10~5_combout ),
	.cin(gnd),
	.combout(Selector101),
	.cout());
// synopsys translate_off
defparam \Selector10~6 .lut_mask = 16'hFFF8;
defparam \Selector10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N20
cycloneive_lcell_comb \Selector10~7 (
// Equation(s):
// Selector102 = (Selector8 & ((\ShiftRight0~99_combout ) # ((\Selector0~23_combout  & \ShiftLeft0~103_combout )))) # (!Selector8 & (((\Selector0~23_combout  & \ShiftLeft0~103_combout ))))

	.dataa(Selector8),
	.datab(\ShiftRight0~99_combout ),
	.datac(\Selector0~23_combout ),
	.datad(\ShiftLeft0~103_combout ),
	.cin(gnd),
	.combout(Selector102),
	.cout());
// synopsys translate_off
defparam \Selector10~7 .lut_mask = 16'hF888;
defparam \Selector10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N18
cycloneive_lcell_comb \Selector10~8 (
// Equation(s):
// Selector103 = (Selector102) # ((Selector10) # (Selector101))

	.dataa(gnd),
	.datab(Selector102),
	.datac(Selector10),
	.datad(Selector101),
	.cin(gnd),
	.combout(Selector103),
	.cout());
// synopsys translate_off
defparam \Selector10~8 .lut_mask = 16'hFFFC;
defparam \Selector10~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N8
cycloneive_lcell_comb \Selector2~9 (
// Equation(s):
// Selector2 = (\Selector2~8_combout ) # ((\Selector2~6_combout ) # ((\Add1~58_combout  & \Selector0~14_combout )))

	.dataa(\Selector2~8_combout ),
	.datab(\Add1~58_combout ),
	.datac(\Selector0~14_combout ),
	.datad(\Selector2~6_combout ),
	.cin(gnd),
	.combout(Selector2),
	.cout());
// synopsys translate_off
defparam \Selector2~9 .lut_mask = 16'hFFEA;
defparam \Selector2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N24
cycloneive_lcell_comb \Selector1~24 (
// Equation(s):
// Selector1 = (\Selector1~18_combout ) # ((\Selector1~12_combout ) # ((\Selector1~23_combout ) # (\Selector1~15_combout )))

	.dataa(\Selector1~18_combout ),
	.datab(\Selector1~12_combout ),
	.datac(\Selector1~23_combout ),
	.datad(\Selector1~15_combout ),
	.cin(gnd),
	.combout(Selector1),
	.cout());
// synopsys translate_off
defparam \Selector1~24 .lut_mask = 16'hFFFE;
defparam \Selector1~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N10
cycloneive_lcell_comb \Selector4~10 (
// Equation(s):
// Selector41 = (\Selector4~9_combout ) # ((\Selector4~6_combout ) # ((Selector4 & \ShiftRight0~125_combout )))

	.dataa(Selector4),
	.datab(\ShiftRight0~125_combout ),
	.datac(\Selector4~9_combout ),
	.datad(\Selector4~6_combout ),
	.cin(gnd),
	.combout(Selector41),
	.cout());
// synopsys translate_off
defparam \Selector4~10 .lut_mask = 16'hFFF8;
defparam \Selector4~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N6
cycloneive_lcell_comb \Selector5~7 (
// Equation(s):
// Selector5 = (\Selector5~4_combout ) # ((\Selector5~1_combout ) # ((\Selector4~0_combout  & \Selector5~6_combout )))

	.dataa(\Selector4~0_combout ),
	.datab(\Selector5~4_combout ),
	.datac(\Selector5~6_combout ),
	.datad(\Selector5~1_combout ),
	.cin(gnd),
	.combout(Selector5),
	.cout());
// synopsys translate_off
defparam \Selector5~7 .lut_mask = 16'hFFEC;
defparam \Selector5~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N12
cycloneive_lcell_comb \Selector5~8 (
// Equation(s):
// Selector51 = (Selector5) # ((Selector4 & ShiftRight02))

	.dataa(Selector4),
	.datab(ShiftRight02),
	.datac(gnd),
	.datad(Selector5),
	.cin(gnd),
	.combout(Selector51),
	.cout());
// synopsys translate_off
defparam \Selector5~8 .lut_mask = 16'hFF88;
defparam \Selector5~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N4
cycloneive_lcell_comb \Selector12~8 (
// Equation(s):
// Selector12 = (\Selector12~1_combout ) # ((\Selector12~7_combout ) # ((Selector8 & \ShiftRight0~74_combout )))

	.dataa(Selector8),
	.datab(\Selector12~1_combout ),
	.datac(\Selector12~7_combout ),
	.datad(\ShiftRight0~74_combout ),
	.cin(gnd),
	.combout(Selector12),
	.cout());
// synopsys translate_off
defparam \Selector12~8 .lut_mask = 16'hFEFC;
defparam \Selector12~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N16
cycloneive_lcell_comb \Selector24~9 (
// Equation(s):
// Selector241 = (\Selector0~9_combout  & (!Mux28 & (!Mux272 & !\ShiftRight0~22_combout )))

	.dataa(\Selector0~9_combout ),
	.datab(Mux28),
	.datac(Mux272),
	.datad(\ShiftRight0~22_combout ),
	.cin(gnd),
	.combout(Selector241),
	.cout());
// synopsys translate_off
defparam \Selector24~9 .lut_mask = 16'h0002;
defparam \Selector24~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N20
cycloneive_lcell_comb \Selector24~10 (
// Equation(s):
// Selector242 = (\Selector24~8_combout ) # ((\Selector24~5_combout ) # ((Selector241 & \ShiftLeft0~101_combout )))

	.dataa(\Selector24~8_combout ),
	.datab(Selector241),
	.datac(\Selector24~5_combout ),
	.datad(\ShiftLeft0~101_combout ),
	.cin(gnd),
	.combout(Selector242),
	.cout());
// synopsys translate_off
defparam \Selector24~10 .lut_mask = 16'hFEFA;
defparam \Selector24~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N4
cycloneive_lcell_comb \Selector13~8 (
// Equation(s):
// Selector13 = (\Selector13~1_combout ) # ((\Selector13~7_combout ) # ((Selector8 & ShiftRight03)))

	.dataa(Selector8),
	.datab(\Selector13~1_combout ),
	.datac(\Selector13~7_combout ),
	.datad(ShiftRight03),
	.cin(gnd),
	.combout(Selector13),
	.cout());
// synopsys translate_off
defparam \Selector13~8 .lut_mask = 16'hFEFC;
defparam \Selector13~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N28
cycloneive_lcell_comb \Selector25~8 (
// Equation(s):
// Selector25 = (\Selector25~7_combout ) # ((\Selector25~4_combout ) # ((Selector241 & \ShiftLeft0~74_combout )))

	.dataa(Selector241),
	.datab(\Selector25~7_combout ),
	.datac(\ShiftLeft0~74_combout ),
	.datad(\Selector25~4_combout ),
	.cin(gnd),
	.combout(Selector25),
	.cout());
// synopsys translate_off
defparam \Selector25~8 .lut_mask = 16'hFFEC;
defparam \Selector25~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N26
cycloneive_lcell_comb \Selector14~1 (
// Equation(s):
// Selector14 = (\ShiftLeft0~94_combout  & ((\Selector8~2_combout ) # ((\Selector0~22_combout  & \Selector14~0_combout )))) # (!\ShiftLeft0~94_combout  & (\Selector0~22_combout  & (\Selector14~0_combout )))

	.dataa(\ShiftLeft0~94_combout ),
	.datab(\Selector0~22_combout ),
	.datac(\Selector14~0_combout ),
	.datad(\Selector8~2_combout ),
	.cin(gnd),
	.combout(Selector14),
	.cout());
// synopsys translate_off
defparam \Selector14~1 .lut_mask = 16'hEAC0;
defparam \Selector14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N30
cycloneive_lcell_comb \Selector14~6 (
// Equation(s):
// Selector141 = (\Selector14~5_combout ) # ((\Selector14~2_combout ) # ((\Selector0~17_combout  & Mux14)))

	.dataa(\Selector0~17_combout ),
	.datab(Mux14),
	.datac(\Selector14~5_combout ),
	.datad(\Selector14~2_combout ),
	.cin(gnd),
	.combout(Selector141),
	.cout());
// synopsys translate_off
defparam \Selector14~6 .lut_mask = 16'hFFF8;
defparam \Selector14~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N26
cycloneive_lcell_comb \Selector14~7 (
// Equation(s):
// Selector142 = (\Selector0~23_combout  & ((\ShiftLeft0~95_combout ) # ((Selector8 & \ShiftRight0~112_combout )))) # (!\Selector0~23_combout  & (Selector8 & ((\ShiftRight0~112_combout ))))

	.dataa(\Selector0~23_combout ),
	.datab(Selector8),
	.datac(\ShiftLeft0~95_combout ),
	.datad(\ShiftRight0~112_combout ),
	.cin(gnd),
	.combout(Selector142),
	.cout());
// synopsys translate_off
defparam \Selector14~7 .lut_mask = 16'hECA0;
defparam \Selector14~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N8
cycloneive_lcell_comb \Selector14~8 (
// Equation(s):
// Selector143 = (Selector14) # ((Selector141) # (Selector142))

	.dataa(gnd),
	.datab(Selector14),
	.datac(Selector141),
	.datad(Selector142),
	.cin(gnd),
	.combout(Selector143),
	.cout());
// synopsys translate_off
defparam \Selector14~8 .lut_mask = 16'hFFFC;
defparam \Selector14~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N16
cycloneive_lcell_comb \Selector27~8 (
// Equation(s):
// Selector27 = (\Selector27~7_combout ) # ((\Selector27~4_combout ) # ((\ShiftLeft0~102_combout  & Selector241)))

	.dataa(\ShiftLeft0~102_combout ),
	.datab(\Selector27~7_combout ),
	.datac(\Selector27~4_combout ),
	.datad(Selector241),
	.cin(gnd),
	.combout(Selector27),
	.cout());
// synopsys translate_off
defparam \Selector27~8 .lut_mask = 16'hFEFC;
defparam \Selector27~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N16
cycloneive_lcell_comb \Selector16~11 (
// Equation(s):
// Selector16 = (\Selector16~6_combout ) # ((\Selector16~10_combout ) # ((\Selector16~1_combout  & \ShiftLeft0~96_combout )))

	.dataa(\Selector16~1_combout ),
	.datab(\ShiftLeft0~96_combout ),
	.datac(\Selector16~6_combout ),
	.datad(\Selector16~10_combout ),
	.cin(gnd),
	.combout(Selector16),
	.cout());
// synopsys translate_off
defparam \Selector16~11 .lut_mask = 16'hFFF8;
defparam \Selector16~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N22
cycloneive_lcell_comb \Selector18~8 (
// Equation(s):
// Selector18 = (\Selector18~1_combout ) # ((\Selector18~7_combout ) # ((\Selector16~1_combout  & \ShiftLeft0~97_combout )))

	.dataa(\Selector16~1_combout ),
	.datab(\Selector18~1_combout ),
	.datac(\Selector18~7_combout ),
	.datad(\ShiftLeft0~97_combout ),
	.cin(gnd),
	.combout(Selector18),
	.cout());
// synopsys translate_off
defparam \Selector18~8 .lut_mask = 16'hFEFC;
defparam \Selector18~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N22
cycloneive_lcell_comb \Selector17~8 (
// Equation(s):
// Selector17 = (\Selector17~1_combout ) # ((\Selector17~7_combout ) # ((\Selector16~1_combout  & \ShiftLeft0~98_combout )))

	.dataa(\Selector16~1_combout ),
	.datab(\ShiftLeft0~98_combout ),
	.datac(\Selector17~1_combout ),
	.datad(\Selector17~7_combout ),
	.cin(gnd),
	.combout(Selector17),
	.cout());
// synopsys translate_off
defparam \Selector17~8 .lut_mask = 16'hFFF8;
defparam \Selector17~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N4
cycloneive_lcell_comb \Selector6~7 (
// Equation(s):
// Selector6 = (\Selector6~2_combout ) # ((\Selector6~6_combout ) # ((\Selector4~0_combout  & \Selector6~1_combout )))

	.dataa(\Selector6~2_combout ),
	.datab(\Selector4~0_combout ),
	.datac(\Selector6~6_combout ),
	.datad(\Selector6~1_combout ),
	.cin(gnd),
	.combout(Selector6),
	.cout());
// synopsys translate_off
defparam \Selector6~7 .lut_mask = 16'hFEFA;
defparam \Selector6~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N28
cycloneive_lcell_comb \Selector26~7 (
// Equation(s):
// Selector26 = (\Selector26~1_combout ) # ((\Selector26~4_combout ) # ((Selector24 & \Selector26~6_combout )))

	.dataa(Selector24),
	.datab(\Selector26~1_combout ),
	.datac(\Selector26~4_combout ),
	.datad(\Selector26~6_combout ),
	.cin(gnd),
	.combout(Selector26),
	.cout());
// synopsys translate_off
defparam \Selector26~7 .lut_mask = 16'hFEFC;
defparam \Selector26~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N2
cycloneive_lcell_comb \Selector26~8 (
// Equation(s):
// Selector261 = (Selector26) # ((Selector241 & ShiftLeft0))

	.dataa(gnd),
	.datab(Selector241),
	.datac(ShiftLeft0),
	.datad(Selector26),
	.cin(gnd),
	.combout(Selector261),
	.cout());
// synopsys translate_off
defparam \Selector26~8 .lut_mask = 16'hFFC0;
defparam \Selector26~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N8
cycloneive_lcell_comb \Selector19~8 (
// Equation(s):
// Selector19 = (\Selector19~1_combout ) # ((\Selector19~7_combout ) # ((\ShiftLeft0~48_combout  & \Selector16~1_combout )))

	.dataa(\ShiftLeft0~48_combout ),
	.datab(\Selector16~1_combout ),
	.datac(\Selector19~1_combout ),
	.datad(\Selector19~7_combout ),
	.cin(gnd),
	.combout(Selector19),
	.cout());
// synopsys translate_off
defparam \Selector19~8 .lut_mask = 16'hFFF8;
defparam \Selector19~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N18
cycloneive_lcell_comb \Selector20~2 (
// Equation(s):
// Selector20 = (\Selector20~1_combout  & ((\ShiftRight0~125_combout ) # ((\Selector0~35_combout  & \Selector20~0_combout )))) # (!\Selector20~1_combout  & (((\Selector0~35_combout  & \Selector20~0_combout ))))

	.dataa(\Selector20~1_combout ),
	.datab(\ShiftRight0~125_combout ),
	.datac(\Selector0~35_combout ),
	.datad(\Selector20~0_combout ),
	.cin(gnd),
	.combout(Selector20),
	.cout());
// synopsys translate_off
defparam \Selector20~2 .lut_mask = 16'hF888;
defparam \Selector20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N24
cycloneive_lcell_comb \Selector20~7 (
// Equation(s):
// Selector201 = (\Selector20~3_combout ) # ((\Selector20~6_combout ) # ((\Selector0~17_combout  & Mux20)))

	.dataa(\Selector20~3_combout ),
	.datab(\Selector0~17_combout ),
	.datac(\Selector20~6_combout ),
	.datad(Mux20),
	.cin(gnd),
	.combout(Selector201),
	.cout());
// synopsys translate_off
defparam \Selector20~7 .lut_mask = 16'hFEFA;
defparam \Selector20~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N30
cycloneive_lcell_comb \Selector20~8 (
// Equation(s):
// Selector202 = (\Selector16~1_combout  & ((\ShiftLeft0~90_combout ) # ((\ShiftRight0~64_combout  & \Selector16~9_combout )))) # (!\Selector16~1_combout  & (\ShiftRight0~64_combout  & (\Selector16~9_combout )))

	.dataa(\Selector16~1_combout ),
	.datab(\ShiftRight0~64_combout ),
	.datac(\Selector16~9_combout ),
	.datad(\ShiftLeft0~90_combout ),
	.cin(gnd),
	.combout(Selector202),
	.cout());
// synopsys translate_off
defparam \Selector20~8 .lut_mask = 16'hEAC0;
defparam \Selector20~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N0
cycloneive_lcell_comb \Selector21~1 (
// Equation(s):
// Selector21 = (ShiftRight02 & ((\Selector20~1_combout ) # ((\Selector21~0_combout  & \Selector0~35_combout )))) # (!ShiftRight02 & (((\Selector21~0_combout  & \Selector0~35_combout ))))

	.dataa(ShiftRight02),
	.datab(\Selector20~1_combout ),
	.datac(\Selector21~0_combout ),
	.datad(\Selector0~35_combout ),
	.cin(gnd),
	.combout(Selector21),
	.cout());
// synopsys translate_off
defparam \Selector21~1 .lut_mask = 16'hF888;
defparam \Selector21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N20
cycloneive_lcell_comb \Selector21~6 (
// Equation(s):
// Selector211 = (\Selector21~5_combout ) # ((\Selector21~2_combout ) # ((Mux21 & \Selector0~17_combout )))

	.dataa(Mux21),
	.datab(\Selector21~5_combout ),
	.datac(\Selector0~17_combout ),
	.datad(\Selector21~2_combout ),
	.cin(gnd),
	.combout(Selector211),
	.cout());
// synopsys translate_off
defparam \Selector21~6 .lut_mask = 16'hFFEC;
defparam \Selector21~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N2
cycloneive_lcell_comb \Selector21~7 (
// Equation(s):
// Selector212 = (\Selector16~9_combout  & ((\ShiftRight0~81_combout ) # ((\Selector16~1_combout  & \ShiftLeft0~93_combout )))) # (!\Selector16~9_combout  & (\Selector16~1_combout  & ((\ShiftLeft0~93_combout ))))

	.dataa(\Selector16~9_combout ),
	.datab(\Selector16~1_combout ),
	.datac(\ShiftRight0~81_combout ),
	.datad(\ShiftLeft0~93_combout ),
	.cin(gnd),
	.combout(Selector212),
	.cout());
// synopsys translate_off
defparam \Selector21~7 .lut_mask = 16'hECA0;
defparam \Selector21~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N30
cycloneive_lcell_comb \Selector21~8 (
// Equation(s):
// Selector213 = (Selector21) # ((Selector212) # (Selector211))

	.dataa(Selector21),
	.datab(gnd),
	.datac(Selector212),
	.datad(Selector211),
	.cin(gnd),
	.combout(Selector213),
	.cout());
// synopsys translate_off
defparam \Selector21~8 .lut_mask = 16'hFFFA;
defparam \Selector21~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N8
cycloneive_lcell_comb \Selector8~3 (
// Equation(s):
// Selector81 = (\Selector8~1_combout  & ((\Selector0~22_combout ) # ((\ShiftLeft0~101_combout  & \Selector8~2_combout )))) # (!\Selector8~1_combout  & (\ShiftLeft0~101_combout  & ((\Selector8~2_combout ))))

	.dataa(\Selector8~1_combout ),
	.datab(\ShiftLeft0~101_combout ),
	.datac(\Selector0~22_combout ),
	.datad(\Selector8~2_combout ),
	.cin(gnd),
	.combout(Selector81),
	.cout());
// synopsys translate_off
defparam \Selector8~3 .lut_mask = 16'hECA0;
defparam \Selector8~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N12
cycloneive_lcell_comb \Selector8~8 (
// Equation(s):
// Selector82 = (\Selector8~7_combout ) # ((\Selector8~4_combout ) # ((Mux8 & \Selector0~17_combout )))

	.dataa(Mux8),
	.datab(\Selector8~7_combout ),
	.datac(\Selector0~17_combout ),
	.datad(\Selector8~4_combout ),
	.cin(gnd),
	.combout(Selector82),
	.cout());
// synopsys translate_off
defparam \Selector8~8 .lut_mask = 16'hFFEC;
defparam \Selector8~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N28
cycloneive_lcell_comb \Selector8~9 (
// Equation(s):
// Selector83 = (\Selector0~23_combout  & ((\Selector0~36_combout ) # ((Selector8 & \ShiftRight0~103_combout )))) # (!\Selector0~23_combout  & (Selector8 & ((\ShiftRight0~103_combout ))))

	.dataa(\Selector0~23_combout ),
	.datab(Selector8),
	.datac(\Selector0~36_combout ),
	.datad(\ShiftRight0~103_combout ),
	.cin(gnd),
	.combout(Selector83),
	.cout());
// synopsys translate_off
defparam \Selector8~9 .lut_mask = 16'hECA0;
defparam \Selector8~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N26
cycloneive_lcell_comb \Selector8~10 (
// Equation(s):
// Selector84 = (Selector81) # ((Selector83) # (Selector82))

	.dataa(gnd),
	.datab(Selector81),
	.datac(Selector83),
	.datad(Selector82),
	.cin(gnd),
	.combout(Selector84),
	.cout());
// synopsys translate_off
defparam \Selector8~10 .lut_mask = 16'hFFFC;
defparam \Selector8~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N28
cycloneive_lcell_comb \Selector9~1 (
// Equation(s):
// Selector9 = (\ShiftLeft0~74_combout  & ((\Selector8~2_combout ) # ((\Selector9~0_combout  & \Selector0~22_combout )))) # (!\ShiftLeft0~74_combout  & (((\Selector9~0_combout  & \Selector0~22_combout ))))

	.dataa(\ShiftLeft0~74_combout ),
	.datab(\Selector8~2_combout ),
	.datac(\Selector9~0_combout ),
	.datad(\Selector0~22_combout ),
	.cin(gnd),
	.combout(Selector9),
	.cout());
// synopsys translate_off
defparam \Selector9~1 .lut_mask = 16'hF888;
defparam \Selector9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N8
cycloneive_lcell_comb \Selector9~6 (
// Equation(s):
// Selector91 = (\Selector9~5_combout ) # ((\Selector9~2_combout ) # ((\Selector0~17_combout  & Mux9)))

	.dataa(\Selector9~5_combout ),
	.datab(\Selector0~17_combout ),
	.datac(Mux9),
	.datad(\Selector9~2_combout ),
	.cin(gnd),
	.combout(Selector91),
	.cout());
// synopsys translate_off
defparam \Selector9~6 .lut_mask = 16'hFFEA;
defparam \Selector9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N22
cycloneive_lcell_comb \Selector9~7 (
// Equation(s):
// Selector92 = (\Selector1~26_combout  & ((\Selector0~23_combout ) # ((Selector8 & \ShiftRight0~108_combout )))) # (!\Selector1~26_combout  & (Selector8 & ((\ShiftRight0~108_combout ))))

	.dataa(\Selector1~26_combout ),
	.datab(Selector8),
	.datac(\Selector0~23_combout ),
	.datad(\ShiftRight0~108_combout ),
	.cin(gnd),
	.combout(Selector92),
	.cout());
// synopsys translate_off
defparam \Selector9~7 .lut_mask = 16'hECA0;
defparam \Selector9~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N10
cycloneive_lcell_comb \Selector9~8 (
// Equation(s):
// Selector93 = (Selector9) # ((Selector91) # (Selector92))

	.dataa(Selector9),
	.datab(gnd),
	.datac(Selector91),
	.datad(Selector92),
	.cin(gnd),
	.combout(Selector93),
	.cout());
// synopsys translate_off
defparam \Selector9~8 .lut_mask = 16'hFFFA;
defparam \Selector9~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N28
cycloneive_lcell_comb \Selector22~9 (
// Equation(s):
// Selector221 = (\Selector22~2_combout ) # ((\Selector22~7_combout ) # ((\Selector22~4_combout ) # (\Selector22~8_combout )))

	.dataa(\Selector22~2_combout ),
	.datab(\Selector22~7_combout ),
	.datac(\Selector22~4_combout ),
	.datad(\Selector22~8_combout ),
	.cin(gnd),
	.combout(Selector221),
	.cout());
// synopsys translate_off
defparam \Selector22~9 .lut_mask = 16'hFFFE;
defparam \Selector22~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N10
cycloneive_lcell_comb \Selector30~14 (
// Equation(s):
// Selector30 = (\Selector30~9_combout ) # ((Selector24 & (!Mux272 & \Selector30~13_combout )))

	.dataa(Selector24),
	.datab(Mux272),
	.datac(\Selector30~9_combout ),
	.datad(\Selector30~13_combout ),
	.cin(gnd),
	.combout(Selector30),
	.cout());
// synopsys translate_off
defparam \Selector30~14 .lut_mask = 16'hF2F0;
defparam \Selector30~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N12
cycloneive_lcell_comb \Selector23~3 (
// Equation(s):
// Selector23 = (\ShiftRight0~121_combout  & ((\Selector16~9_combout ) # ((\Selector20~1_combout  & \ShiftRight0~30_combout )))) # (!\ShiftRight0~121_combout  & (\Selector20~1_combout  & ((\ShiftRight0~30_combout ))))

	.dataa(\ShiftRight0~121_combout ),
	.datab(\Selector20~1_combout ),
	.datac(\Selector16~9_combout ),
	.datad(\ShiftRight0~30_combout ),
	.cin(gnd),
	.combout(Selector23),
	.cout());
// synopsys translate_off
defparam \Selector23~3 .lut_mask = 16'hECA0;
defparam \Selector23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N26
cycloneive_lcell_comb \Selector23~4 (
// Equation(s):
// Selector231 = (\Selector0~35_combout  & \Selector23~2_combout )

	.dataa(gnd),
	.datab(\Selector0~35_combout ),
	.datac(gnd),
	.datad(\Selector23~2_combout ),
	.cin(gnd),
	.combout(Selector231),
	.cout());
// synopsys translate_off
defparam \Selector23~4 .lut_mask = 16'hCC00;
defparam \Selector23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N16
cycloneive_lcell_comb \Selector23~10 (
// Equation(s):
// Selector232 = (\Selector23~9_combout ) # ((\ShiftLeft0~51_combout  & \Selector16~1_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~51_combout ),
	.datac(\Selector23~9_combout ),
	.datad(\Selector16~1_combout ),
	.cin(gnd),
	.combout(Selector232),
	.cout());
// synopsys translate_off
defparam \Selector23~10 .lut_mask = 16'hFCF0;
defparam \Selector23~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N6
cycloneive_lcell_comb \Equal0~11 (
// Equation(s):
// Equal0 = (\Equal0~3_combout  & (\Equal0~10_combout  & (\Equal0~8_combout  & \Equal0~9_combout )))

	.dataa(\Equal0~3_combout ),
	.datab(\Equal0~10_combout ),
	.datac(\Equal0~8_combout ),
	.datad(\Equal0~9_combout ),
	.cin(gnd),
	.combout(Equal0),
	.cout());
// synopsys translate_off
defparam \Equal0~11 .lut_mask = 16'h8000;
defparam \Equal0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N14
cycloneive_lcell_comb \Selector20~9 (
// Equation(s):
// Selector203 = (Selector202) # ((Selector20) # (Selector201))

	.dataa(Selector202),
	.datab(Selector20),
	.datac(gnd),
	.datad(Selector201),
	.cin(gnd),
	.combout(Selector203),
	.cout());
// synopsys translate_off
defparam \Selector20~9 .lut_mask = 16'hFFEE;
defparam \Selector20~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N10
cycloneive_lcell_comb \Selector31~12 (
// Equation(s):
// Selector311 = (Selector31) # ((!\ShiftRight0~22_combout  & (\Selector0~13_combout  & ShiftRight0)))

	.dataa(\ShiftRight0~22_combout ),
	.datab(\Selector0~13_combout ),
	.datac(ShiftRight0),
	.datad(Selector31),
	.cin(gnd),
	.combout(Selector311),
	.cout());
// synopsys translate_off
defparam \Selector31~12 .lut_mask = 16'hFF40;
defparam \Selector31~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N10
cycloneive_lcell_comb \Selector23~11 (
// Equation(s):
// Selector233 = (Selector23) # ((Selector232) # ((\Selector23~2_combout  & \Selector0~35_combout )))

	.dataa(\Selector23~2_combout ),
	.datab(\Selector0~35_combout ),
	.datac(Selector23),
	.datad(Selector232),
	.cin(gnd),
	.combout(Selector233),
	.cout());
// synopsys translate_off
defparam \Selector23~11 .lut_mask = 16'hFFF8;
defparam \Selector23~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N14
cycloneive_lcell_comb \Selector0~4 (
// Equation(s):
// \Selector0~4_combout  = (cuifALUOP_0 & (cuifALUOP_3 & (cuifALUOP_1 & !cuifALUOP_2)))

	.dataa(cuifALUOP_0),
	.datab(cuifALUOP_3),
	.datac(cuifALUOP_1),
	.datad(cuifALUOP_2),
	.cin(gnd),
	.combout(\Selector0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~4 .lut_mask = 16'h0080;
defparam \Selector0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N10
cycloneive_lcell_comb \Selector0~5 (
// Equation(s):
// \Selector0~5_combout  = (cuifALUOP_0 & (!cuifALUOP_1 & (!cuifALUOP_3 & cuifALUOP_2)))

	.dataa(cuifALUOP_0),
	.datab(cuifALUOP_1),
	.datac(cuifALUOP_3),
	.datad(cuifALUOP_2),
	.cin(gnd),
	.combout(\Selector0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~5 .lut_mask = 16'h0200;
defparam \Selector0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N0
cycloneive_lcell_comb \Selector0~6 (
// Equation(s):
// \Selector0~6_combout  = (!cuifALUOP_1 & (!cuifALUOP_3 & (!cuifALUOP_0 & cuifALUOP_2)))

	.dataa(cuifALUOP_1),
	.datab(cuifALUOP_3),
	.datac(cuifALUOP_0),
	.datad(cuifALUOP_2),
	.cin(gnd),
	.combout(\Selector0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~6 .lut_mask = 16'h0100;
defparam \Selector0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N2
cycloneive_lcell_comb \Selector31~4 (
// Equation(s):
// \Selector31~4_combout  = (\Selector0~5_combout ) # ((Mux312 & \Selector0~6_combout ))

	.dataa(Mux312),
	.datab(\Selector0~5_combout ),
	.datac(gnd),
	.datad(\Selector0~6_combout ),
	.cin(gnd),
	.combout(\Selector31~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~4 .lut_mask = 16'hEECC;
defparam \Selector31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N0
cycloneive_lcell_comb \Add1~0 (
// Equation(s):
// \Add1~0_combout  = (\portB~65_combout  & (Mux312 $ (VCC))) # (!\portB~65_combout  & ((Mux312) # (GND)))
// \Add1~1  = CARRY((Mux312) # (!\portB~65_combout ))

	.dataa(portB31),
	.datab(Mux312),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h66DD;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N16
cycloneive_lcell_comb \Selector0~8 (
// Equation(s):
// \Selector0~8_combout  = (cuifALUOP_1 & (!cuifALUOP_3 & (cuifALUOP_0 & !cuifALUOP_2)))

	.dataa(cuifALUOP_1),
	.datab(cuifALUOP_3),
	.datac(cuifALUOP_0),
	.datad(cuifALUOP_2),
	.cin(gnd),
	.combout(\Selector0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~8 .lut_mask = 16'h0020;
defparam \Selector0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N0
cycloneive_lcell_comb \ShiftRight0~23 (
// Equation(s):
// \ShiftRight0~23_combout  = (Mux312) # ((Mux292) # ((Mux28) # (Mux302)))

	.dataa(Mux312),
	.datab(Mux292),
	.datac(Mux28),
	.datad(Mux302),
	.cin(gnd),
	.combout(\ShiftRight0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~23 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N20
cycloneive_lcell_comb \Selector0~9 (
// Equation(s):
// \Selector0~9_combout  = (!cuifALUOP_2 & (!cuifALUOP_1 & (!cuifALUOP_0 & !cuifALUOP_3)))

	.dataa(cuifALUOP_2),
	.datab(cuifALUOP_1),
	.datac(cuifALUOP_0),
	.datad(cuifALUOP_3),
	.cin(gnd),
	.combout(\Selector0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~9 .lut_mask = 16'h0001;
defparam \Selector0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N28
cycloneive_lcell_comb \ShiftRight0~20 (
// Equation(s):
// \ShiftRight0~20_combout  = (Mux21) # ((Mux20) # ((Mux22) # (Mux23)))

	.dataa(Mux21),
	.datab(Mux20),
	.datac(Mux22),
	.datad(Mux23),
	.cin(gnd),
	.combout(\ShiftRight0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~20 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N18
cycloneive_lcell_comb \ShiftRight0~14 (
// Equation(s):
// \ShiftRight0~14_combout  = (Mux1) # ((Mux0) # ((Mux3) # (Mux2)))

	.dataa(Mux1),
	.datab(Mux0),
	.datac(Mux3),
	.datad(Mux2),
	.cin(gnd),
	.combout(\ShiftRight0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~14 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N4
cycloneive_lcell_comb \ShiftRight0~17 (
// Equation(s):
// \ShiftRight0~17_combout  = (Mux15) # ((Mux13) # ((Mux14) # (Mux12)))

	.dataa(Mux15),
	.datab(Mux13),
	.datac(Mux14),
	.datad(Mux12),
	.cin(gnd),
	.combout(\ShiftRight0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~17 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N14
cycloneive_lcell_comb \ShiftRight0~16 (
// Equation(s):
// \ShiftRight0~16_combout  = (Mux8) # ((Mux10) # ((Mux9) # (Mux11)))

	.dataa(Mux8),
	.datab(Mux10),
	.datac(Mux9),
	.datad(Mux11),
	.cin(gnd),
	.combout(\ShiftRight0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~16 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N26
cycloneive_lcell_comb \ShiftRight0~18 (
// Equation(s):
// \ShiftRight0~18_combout  = (\ShiftRight0~15_combout ) # ((\ShiftRight0~14_combout ) # ((\ShiftRight0~17_combout ) # (\ShiftRight0~16_combout )))

	.dataa(\ShiftRight0~15_combout ),
	.datab(\ShiftRight0~14_combout ),
	.datac(\ShiftRight0~17_combout ),
	.datad(\ShiftRight0~16_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~18 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N2
cycloneive_lcell_comb \ShiftRight0~19 (
// Equation(s):
// \ShiftRight0~19_combout  = (Mux19) # ((Mux16) # ((Mux18) # (Mux17)))

	.dataa(Mux19),
	.datab(Mux16),
	.datac(Mux18),
	.datad(Mux17),
	.cin(gnd),
	.combout(\ShiftRight0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~19 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N24
cycloneive_lcell_comb \ShiftRight0~22 (
// Equation(s):
// \ShiftRight0~22_combout  = (\ShiftRight0~21_combout ) # ((\ShiftRight0~20_combout ) # ((\ShiftRight0~18_combout ) # (\ShiftRight0~19_combout )))

	.dataa(\ShiftRight0~21_combout ),
	.datab(\ShiftRight0~20_combout ),
	.datac(\ShiftRight0~18_combout ),
	.datad(\ShiftRight0~19_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~22 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N0
cycloneive_lcell_comb \Selector31~11 (
// Equation(s):
// \Selector31~11_combout  = (!Mux272 & (!\ShiftRight0~23_combout  & (\Selector0~9_combout  & !\ShiftRight0~22_combout )))

	.dataa(Mux272),
	.datab(\ShiftRight0~23_combout ),
	.datac(\Selector0~9_combout ),
	.datad(\ShiftRight0~22_combout ),
	.cin(gnd),
	.combout(\Selector31~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~11 .lut_mask = 16'h0010;
defparam \Selector31~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N14
cycloneive_lcell_comb \Selector31~6 (
// Equation(s):
// \Selector31~6_combout  = (\portB~65_combout  & ((\Selector31~11_combout ) # ((\Add1~0_combout  & \Selector0~8_combout )))) # (!\portB~65_combout  & (\Add1~0_combout  & (\Selector0~8_combout )))

	.dataa(portB31),
	.datab(\Add1~0_combout ),
	.datac(\Selector0~8_combout ),
	.datad(\Selector31~11_combout ),
	.cin(gnd),
	.combout(\Selector31~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~6 .lut_mask = 16'hEAC0;
defparam \Selector31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N24
cycloneive_lcell_comb \Selector31~5 (
// Equation(s):
// \Selector31~5_combout  = (Mux312 & (((\Selector0~5_combout )))) # (!Mux312 & (\Selector0~7_combout  & ((!\portB~65_combout ))))

	.dataa(\Selector0~7_combout ),
	.datab(\Selector0~5_combout ),
	.datac(portB31),
	.datad(Mux312),
	.cin(gnd),
	.combout(\Selector31~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~5 .lut_mask = 16'hCC0A;
defparam \Selector31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N16
cycloneive_lcell_comb \Selector31~7 (
// Equation(s):
// \Selector31~7_combout  = (\Selector31~6_combout ) # ((\Selector31~5_combout ) # ((\portB~65_combout  & \Selector31~4_combout )))

	.dataa(portB31),
	.datab(\Selector31~4_combout ),
	.datac(\Selector31~6_combout ),
	.datad(\Selector31~5_combout ),
	.cin(gnd),
	.combout(\Selector31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~7 .lut_mask = 16'hFFF8;
defparam \Selector31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N28
cycloneive_lcell_comb \Selector0~12 (
// Equation(s):
// \Selector0~12_combout  = (cuifALUOP_1 & (!cuifALUOP_2 & (!cuifALUOP_0 & cuifALUOP_3)))

	.dataa(cuifALUOP_1),
	.datab(cuifALUOP_2),
	.datac(cuifALUOP_0),
	.datad(cuifALUOP_3),
	.cin(gnd),
	.combout(\Selector0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~12 .lut_mask = 16'h0200;
defparam \Selector0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N0
cycloneive_lcell_comb \Add0~0 (
// Equation(s):
// \Add0~0_combout  = (\portB~65_combout  & (Mux312 $ (VCC))) # (!\portB~65_combout  & (Mux312 & VCC))
// \Add0~1  = CARRY((\portB~65_combout  & Mux312))

	.dataa(portB31),
	.datab(Mux312),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
// synopsys translate_off
defparam \Add0~0 .lut_mask = 16'h6688;
defparam \Add0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N8
cycloneive_lcell_comb \Selector0~11 (
// Equation(s):
// \Selector0~11_combout  = (cuifALUOP_2 & (!cuifALUOP_0 & (!cuifALUOP_3 & cuifALUOP_1)))

	.dataa(cuifALUOP_2),
	.datab(cuifALUOP_0),
	.datac(cuifALUOP_3),
	.datad(cuifALUOP_1),
	.cin(gnd),
	.combout(\Selector0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~11 .lut_mask = 16'h0200;
defparam \Selector0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N0
cycloneive_lcell_comb \Selector31~8 (
// Equation(s):
// \Selector31~8_combout  = (\Add0~0_combout  & ((\Selector0~10_combout ) # (\Selector0~11_combout )))

	.dataa(\Selector0~10_combout ),
	.datab(gnd),
	.datac(\Add0~0_combout ),
	.datad(\Selector0~11_combout ),
	.cin(gnd),
	.combout(\Selector31~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~8 .lut_mask = 16'hF0A0;
defparam \Selector31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N0
cycloneive_lcell_comb \LessThan0~1 (
// Equation(s):
// \LessThan0~1_cout  = CARRY((!Mux312 & \portB~65_combout ))

	.dataa(Mux312),
	.datab(portB31),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan0~1_cout ));
// synopsys translate_off
defparam \LessThan0~1 .lut_mask = 16'h0044;
defparam \LessThan0~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N2
cycloneive_lcell_comb \LessThan0~3 (
// Equation(s):
// \LessThan0~3_cout  = CARRY((Mux302 & ((!\LessThan0~1_cout ) # (!\portB~63_combout ))) # (!Mux302 & (!\portB~63_combout  & !\LessThan0~1_cout )))

	.dataa(Mux302),
	.datab(portB30),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~1_cout ),
	.combout(),
	.cout(\LessThan0~3_cout ));
// synopsys translate_off
defparam \LessThan0~3 .lut_mask = 16'h002B;
defparam \LessThan0~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N4
cycloneive_lcell_comb \LessThan0~5 (
// Equation(s):
// \LessThan0~5_cout  = CARRY((\portB~61_combout  & ((!\LessThan0~3_cout ) # (!Mux292))) # (!\portB~61_combout  & (!Mux292 & !\LessThan0~3_cout )))

	.dataa(portB29),
	.datab(Mux292),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~3_cout ),
	.combout(),
	.cout(\LessThan0~5_cout ));
// synopsys translate_off
defparam \LessThan0~5 .lut_mask = 16'h002B;
defparam \LessThan0~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N6
cycloneive_lcell_comb \LessThan0~7 (
// Equation(s):
// \LessThan0~7_cout  = CARRY((Mux28 & ((!\LessThan0~5_cout ) # (!\portB~59_combout ))) # (!Mux28 & (!\portB~59_combout  & !\LessThan0~5_cout )))

	.dataa(Mux28),
	.datab(portB28),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~5_cout ),
	.combout(),
	.cout(\LessThan0~7_cout ));
// synopsys translate_off
defparam \LessThan0~7 .lut_mask = 16'h002B;
defparam \LessThan0~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N8
cycloneive_lcell_comb \LessThan0~9 (
// Equation(s):
// \LessThan0~9_cout  = CARRY((Mux272 & (\portB~57_combout  & !\LessThan0~7_cout )) # (!Mux272 & ((\portB~57_combout ) # (!\LessThan0~7_cout ))))

	.dataa(Mux272),
	.datab(portB27),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~7_cout ),
	.combout(),
	.cout(\LessThan0~9_cout ));
// synopsys translate_off
defparam \LessThan0~9 .lut_mask = 16'h004D;
defparam \LessThan0~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N10
cycloneive_lcell_comb \LessThan0~11 (
// Equation(s):
// \LessThan0~11_cout  = CARRY((Mux26 & ((!\LessThan0~9_cout ) # (!\portB~55_combout ))) # (!Mux26 & (!\portB~55_combout  & !\LessThan0~9_cout )))

	.dataa(Mux26),
	.datab(portB26),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~9_cout ),
	.combout(),
	.cout(\LessThan0~11_cout ));
// synopsys translate_off
defparam \LessThan0~11 .lut_mask = 16'h002B;
defparam \LessThan0~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N12
cycloneive_lcell_comb \LessThan0~13 (
// Equation(s):
// \LessThan0~13_cout  = CARRY((Mux252 & (\portB~53_combout  & !\LessThan0~11_cout )) # (!Mux252 & ((\portB~53_combout ) # (!\LessThan0~11_cout ))))

	.dataa(Mux252),
	.datab(portB25),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~11_cout ),
	.combout(),
	.cout(\LessThan0~13_cout ));
// synopsys translate_off
defparam \LessThan0~13 .lut_mask = 16'h004D;
defparam \LessThan0~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N14
cycloneive_lcell_comb \LessThan0~15 (
// Equation(s):
// \LessThan0~15_cout  = CARRY((Mux242 & ((!\LessThan0~13_cout ) # (!\portB~51_combout ))) # (!Mux242 & (!\portB~51_combout  & !\LessThan0~13_cout )))

	.dataa(Mux242),
	.datab(portB24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~13_cout ),
	.combout(),
	.cout(\LessThan0~15_cout ));
// synopsys translate_off
defparam \LessThan0~15 .lut_mask = 16'h002B;
defparam \LessThan0~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N16
cycloneive_lcell_comb \LessThan0~17 (
// Equation(s):
// \LessThan0~17_cout  = CARRY((\portB~49_combout  & ((!\LessThan0~15_cout ) # (!Mux23))) # (!\portB~49_combout  & (!Mux23 & !\LessThan0~15_cout )))

	.dataa(portB23),
	.datab(Mux23),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~15_cout ),
	.combout(),
	.cout(\LessThan0~17_cout ));
// synopsys translate_off
defparam \LessThan0~17 .lut_mask = 16'h002B;
defparam \LessThan0~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N18
cycloneive_lcell_comb \LessThan0~19 (
// Equation(s):
// \LessThan0~19_cout  = CARRY((Mux22 & ((!\LessThan0~17_cout ) # (!\portB~47_combout ))) # (!Mux22 & (!\portB~47_combout  & !\LessThan0~17_cout )))

	.dataa(Mux22),
	.datab(portB22),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~17_cout ),
	.combout(),
	.cout(\LessThan0~19_cout ));
// synopsys translate_off
defparam \LessThan0~19 .lut_mask = 16'h002B;
defparam \LessThan0~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N20
cycloneive_lcell_comb \LessThan0~21 (
// Equation(s):
// \LessThan0~21_cout  = CARRY((\portB~45_combout  & ((!\LessThan0~19_cout ) # (!Mux21))) # (!\portB~45_combout  & (!Mux21 & !\LessThan0~19_cout )))

	.dataa(portB21),
	.datab(Mux21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~19_cout ),
	.combout(),
	.cout(\LessThan0~21_cout ));
// synopsys translate_off
defparam \LessThan0~21 .lut_mask = 16'h002B;
defparam \LessThan0~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N22
cycloneive_lcell_comb \LessThan0~23 (
// Equation(s):
// \LessThan0~23_cout  = CARRY((\portB~43_combout  & (Mux20 & !\LessThan0~21_cout )) # (!\portB~43_combout  & ((Mux20) # (!\LessThan0~21_cout ))))

	.dataa(portB20),
	.datab(Mux20),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~21_cout ),
	.combout(),
	.cout(\LessThan0~23_cout ));
// synopsys translate_off
defparam \LessThan0~23 .lut_mask = 16'h004D;
defparam \LessThan0~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N24
cycloneive_lcell_comb \LessThan0~25 (
// Equation(s):
// \LessThan0~25_cout  = CARRY((Mux19 & (\portB~41_combout  & !\LessThan0~23_cout )) # (!Mux19 & ((\portB~41_combout ) # (!\LessThan0~23_cout ))))

	.dataa(Mux19),
	.datab(portB19),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~23_cout ),
	.combout(),
	.cout(\LessThan0~25_cout ));
// synopsys translate_off
defparam \LessThan0~25 .lut_mask = 16'h004D;
defparam \LessThan0~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N26
cycloneive_lcell_comb \LessThan0~27 (
// Equation(s):
// \LessThan0~27_cout  = CARRY((Mux18 & ((!\LessThan0~25_cout ) # (!\portB~39_combout ))) # (!Mux18 & (!\portB~39_combout  & !\LessThan0~25_cout )))

	.dataa(Mux18),
	.datab(portB18),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~25_cout ),
	.combout(),
	.cout(\LessThan0~27_cout ));
// synopsys translate_off
defparam \LessThan0~27 .lut_mask = 16'h002B;
defparam \LessThan0~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N28
cycloneive_lcell_comb \LessThan0~29 (
// Equation(s):
// \LessThan0~29_cout  = CARRY((Mux17 & (\portB~37_combout  & !\LessThan0~27_cout )) # (!Mux17 & ((\portB~37_combout ) # (!\LessThan0~27_cout ))))

	.dataa(Mux17),
	.datab(portB17),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~27_cout ),
	.combout(),
	.cout(\LessThan0~29_cout ));
// synopsys translate_off
defparam \LessThan0~29 .lut_mask = 16'h004D;
defparam \LessThan0~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N30
cycloneive_lcell_comb \LessThan0~31 (
// Equation(s):
// \LessThan0~31_cout  = CARRY((\portB~35_combout  & (Mux16 & !\LessThan0~29_cout )) # (!\portB~35_combout  & ((Mux16) # (!\LessThan0~29_cout ))))

	.dataa(portB16),
	.datab(Mux16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~29_cout ),
	.combout(),
	.cout(\LessThan0~31_cout ));
// synopsys translate_off
defparam \LessThan0~31 .lut_mask = 16'h004D;
defparam \LessThan0~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N0
cycloneive_lcell_comb \LessThan0~33 (
// Equation(s):
// \LessThan0~33_cout  = CARRY((\portB~33_combout  & ((!\LessThan0~31_cout ) # (!Mux15))) # (!\portB~33_combout  & (!Mux15 & !\LessThan0~31_cout )))

	.dataa(portB15),
	.datab(Mux15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~31_cout ),
	.combout(),
	.cout(\LessThan0~33_cout ));
// synopsys translate_off
defparam \LessThan0~33 .lut_mask = 16'h002B;
defparam \LessThan0~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N2
cycloneive_lcell_comb \LessThan0~35 (
// Equation(s):
// \LessThan0~35_cout  = CARRY((\portB~31_combout  & (Mux14 & !\LessThan0~33_cout )) # (!\portB~31_combout  & ((Mux14) # (!\LessThan0~33_cout ))))

	.dataa(portB14),
	.datab(Mux14),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~33_cout ),
	.combout(),
	.cout(\LessThan0~35_cout ));
// synopsys translate_off
defparam \LessThan0~35 .lut_mask = 16'h004D;
defparam \LessThan0~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N4
cycloneive_lcell_comb \LessThan0~37 (
// Equation(s):
// \LessThan0~37_cout  = CARRY((Mux13 & (\portB~29_combout  & !\LessThan0~35_cout )) # (!Mux13 & ((\portB~29_combout ) # (!\LessThan0~35_cout ))))

	.dataa(Mux13),
	.datab(portB13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~35_cout ),
	.combout(),
	.cout(\LessThan0~37_cout ));
// synopsys translate_off
defparam \LessThan0~37 .lut_mask = 16'h004D;
defparam \LessThan0~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N6
cycloneive_lcell_comb \LessThan0~39 (
// Equation(s):
// \LessThan0~39_cout  = CARRY((Mux12 & ((!\LessThan0~37_cout ) # (!\portB~27_combout ))) # (!Mux12 & (!\portB~27_combout  & !\LessThan0~37_cout )))

	.dataa(Mux12),
	.datab(portB12),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~37_cout ),
	.combout(),
	.cout(\LessThan0~39_cout ));
// synopsys translate_off
defparam \LessThan0~39 .lut_mask = 16'h002B;
defparam \LessThan0~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N8
cycloneive_lcell_comb \LessThan0~41 (
// Equation(s):
// \LessThan0~41_cout  = CARRY((\portB~25_combout  & ((!\LessThan0~39_cout ) # (!Mux11))) # (!\portB~25_combout  & (!Mux11 & !\LessThan0~39_cout )))

	.dataa(portB11),
	.datab(Mux11),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~39_cout ),
	.combout(),
	.cout(\LessThan0~41_cout ));
// synopsys translate_off
defparam \LessThan0~41 .lut_mask = 16'h002B;
defparam \LessThan0~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N10
cycloneive_lcell_comb \LessThan0~43 (
// Equation(s):
// \LessThan0~43_cout  = CARRY((Mux10 & ((!\LessThan0~41_cout ) # (!\portB~23_combout ))) # (!Mux10 & (!\portB~23_combout  & !\LessThan0~41_cout )))

	.dataa(Mux10),
	.datab(portB10),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~41_cout ),
	.combout(),
	.cout(\LessThan0~43_cout ));
// synopsys translate_off
defparam \LessThan0~43 .lut_mask = 16'h002B;
defparam \LessThan0~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N12
cycloneive_lcell_comb \LessThan0~45 (
// Equation(s):
// \LessThan0~45_cout  = CARRY((\portB~21_combout  & ((!\LessThan0~43_cout ) # (!Mux9))) # (!\portB~21_combout  & (!Mux9 & !\LessThan0~43_cout )))

	.dataa(portB9),
	.datab(Mux9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~43_cout ),
	.combout(),
	.cout(\LessThan0~45_cout ));
// synopsys translate_off
defparam \LessThan0~45 .lut_mask = 16'h002B;
defparam \LessThan0~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N14
cycloneive_lcell_comb \LessThan0~47 (
// Equation(s):
// \LessThan0~47_cout  = CARRY((\portB~19_combout  & (Mux8 & !\LessThan0~45_cout )) # (!\portB~19_combout  & ((Mux8) # (!\LessThan0~45_cout ))))

	.dataa(portB8),
	.datab(Mux8),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~45_cout ),
	.combout(),
	.cout(\LessThan0~47_cout ));
// synopsys translate_off
defparam \LessThan0~47 .lut_mask = 16'h004D;
defparam \LessThan0~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N16
cycloneive_lcell_comb \LessThan0~49 (
// Equation(s):
// \LessThan0~49_cout  = CARRY((\portB~17_combout  & ((!\LessThan0~47_cout ) # (!Mux72))) # (!\portB~17_combout  & (!Mux72 & !\LessThan0~47_cout )))

	.dataa(portB7),
	.datab(Mux72),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~47_cout ),
	.combout(),
	.cout(\LessThan0~49_cout ));
// synopsys translate_off
defparam \LessThan0~49 .lut_mask = 16'h002B;
defparam \LessThan0~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N18
cycloneive_lcell_comb \LessThan0~51 (
// Equation(s):
// \LessThan0~51_cout  = CARRY((\portB~15_combout  & (Mux6 & !\LessThan0~49_cout )) # (!\portB~15_combout  & ((Mux6) # (!\LessThan0~49_cout ))))

	.dataa(portB6),
	.datab(Mux6),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~49_cout ),
	.combout(),
	.cout(\LessThan0~51_cout ));
// synopsys translate_off
defparam \LessThan0~51 .lut_mask = 16'h004D;
defparam \LessThan0~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N20
cycloneive_lcell_comb \LessThan0~53 (
// Equation(s):
// \LessThan0~53_cout  = CARRY((Mux5 & (\portB~13_combout  & !\LessThan0~51_cout )) # (!Mux5 & ((\portB~13_combout ) # (!\LessThan0~51_cout ))))

	.dataa(Mux5),
	.datab(portB5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~51_cout ),
	.combout(),
	.cout(\LessThan0~53_cout ));
// synopsys translate_off
defparam \LessThan0~53 .lut_mask = 16'h004D;
defparam \LessThan0~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N22
cycloneive_lcell_comb \LessThan0~55 (
// Equation(s):
// \LessThan0~55_cout  = CARRY((Mux4 & ((!\LessThan0~53_cout ) # (!\portB~11_combout ))) # (!Mux4 & (!\portB~11_combout  & !\LessThan0~53_cout )))

	.dataa(Mux4),
	.datab(portB4),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~53_cout ),
	.combout(),
	.cout(\LessThan0~55_cout ));
// synopsys translate_off
defparam \LessThan0~55 .lut_mask = 16'h002B;
defparam \LessThan0~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N24
cycloneive_lcell_comb \LessThan0~57 (
// Equation(s):
// \LessThan0~57_cout  = CARRY((Mux3 & (\portB~9_combout  & !\LessThan0~55_cout )) # (!Mux3 & ((\portB~9_combout ) # (!\LessThan0~55_cout ))))

	.dataa(Mux3),
	.datab(portB3),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~55_cout ),
	.combout(),
	.cout(\LessThan0~57_cout ));
// synopsys translate_off
defparam \LessThan0~57 .lut_mask = 16'h004D;
defparam \LessThan0~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N26
cycloneive_lcell_comb \LessThan0~59 (
// Equation(s):
// \LessThan0~59_cout  = CARRY((\portB~7_combout  & (Mux2 & !\LessThan0~57_cout )) # (!\portB~7_combout  & ((Mux2) # (!\LessThan0~57_cout ))))

	.dataa(portB2),
	.datab(Mux2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~57_cout ),
	.combout(),
	.cout(\LessThan0~59_cout ));
// synopsys translate_off
defparam \LessThan0~59 .lut_mask = 16'h004D;
defparam \LessThan0~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N28
cycloneive_lcell_comb \LessThan0~61 (
// Equation(s):
// \LessThan0~61_cout  = CARRY((Mux1 & (\portB~5_combout  & !\LessThan0~59_cout )) # (!Mux1 & ((\portB~5_combout ) # (!\LessThan0~59_cout ))))

	.dataa(Mux1),
	.datab(portB1),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~59_cout ),
	.combout(),
	.cout(\LessThan0~61_cout ));
// synopsys translate_off
defparam \LessThan0~61 .lut_mask = 16'h004D;
defparam \LessThan0~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N30
cycloneive_lcell_comb \LessThan0~62 (
// Equation(s):
// \LessThan0~62_combout  = (\portB~3_combout  & (\LessThan0~61_cout  & Mux0)) # (!\portB~3_combout  & ((\LessThan0~61_cout ) # (Mux0)))

	.dataa(portB),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux0),
	.cin(\LessThan0~61_cout ),
	.combout(\LessThan0~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan0~62 .lut_mask = 16'hF550;
defparam \LessThan0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N22
cycloneive_lcell_comb \Selector31~9 (
// Equation(s):
// \Selector31~9_combout  = (\Selector31~8_combout ) # ((\Selector0~12_combout  & \LessThan0~62_combout ))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector31~8_combout ),
	.datac(gnd),
	.datad(\LessThan0~62_combout ),
	.cin(gnd),
	.combout(\Selector31~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~9 .lut_mask = 16'hEECC;
defparam \Selector31~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N0
cycloneive_lcell_comb \LessThan1~1 (
// Equation(s):
// \LessThan1~1_cout  = CARRY((\portB~65_combout  & !Mux312))

	.dataa(portB31),
	.datab(Mux312),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan1~1_cout ));
// synopsys translate_off
defparam \LessThan1~1 .lut_mask = 16'h0022;
defparam \LessThan1~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N2
cycloneive_lcell_comb \LessThan1~3 (
// Equation(s):
// \LessThan1~3_cout  = CARRY((\portB~63_combout  & (Mux302 & !\LessThan1~1_cout )) # (!\portB~63_combout  & ((Mux302) # (!\LessThan1~1_cout ))))

	.dataa(portB30),
	.datab(Mux302),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~1_cout ),
	.combout(),
	.cout(\LessThan1~3_cout ));
// synopsys translate_off
defparam \LessThan1~3 .lut_mask = 16'h004D;
defparam \LessThan1~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N4
cycloneive_lcell_comb \LessThan1~5 (
// Equation(s):
// \LessThan1~5_cout  = CARRY((Mux292 & (\portB~61_combout  & !\LessThan1~3_cout )) # (!Mux292 & ((\portB~61_combout ) # (!\LessThan1~3_cout ))))

	.dataa(Mux292),
	.datab(portB29),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~3_cout ),
	.combout(),
	.cout(\LessThan1~5_cout ));
// synopsys translate_off
defparam \LessThan1~5 .lut_mask = 16'h004D;
defparam \LessThan1~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N6
cycloneive_lcell_comb \LessThan1~7 (
// Equation(s):
// \LessThan1~7_cout  = CARRY((Mux28 & ((!\LessThan1~5_cout ) # (!\portB~59_combout ))) # (!Mux28 & (!\portB~59_combout  & !\LessThan1~5_cout )))

	.dataa(Mux28),
	.datab(portB28),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~5_cout ),
	.combout(),
	.cout(\LessThan1~7_cout ));
// synopsys translate_off
defparam \LessThan1~7 .lut_mask = 16'h002B;
defparam \LessThan1~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N8
cycloneive_lcell_comb \LessThan1~9 (
// Equation(s):
// \LessThan1~9_cout  = CARRY((Mux272 & (\portB~57_combout  & !\LessThan1~7_cout )) # (!Mux272 & ((\portB~57_combout ) # (!\LessThan1~7_cout ))))

	.dataa(Mux272),
	.datab(portB27),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~7_cout ),
	.combout(),
	.cout(\LessThan1~9_cout ));
// synopsys translate_off
defparam \LessThan1~9 .lut_mask = 16'h004D;
defparam \LessThan1~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N10
cycloneive_lcell_comb \LessThan1~11 (
// Equation(s):
// \LessThan1~11_cout  = CARRY((Mux26 & ((!\LessThan1~9_cout ) # (!\portB~55_combout ))) # (!Mux26 & (!\portB~55_combout  & !\LessThan1~9_cout )))

	.dataa(Mux26),
	.datab(portB26),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~9_cout ),
	.combout(),
	.cout(\LessThan1~11_cout ));
// synopsys translate_off
defparam \LessThan1~11 .lut_mask = 16'h002B;
defparam \LessThan1~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N12
cycloneive_lcell_comb \LessThan1~13 (
// Equation(s):
// \LessThan1~13_cout  = CARRY((Mux252 & (\portB~53_combout  & !\LessThan1~11_cout )) # (!Mux252 & ((\portB~53_combout ) # (!\LessThan1~11_cout ))))

	.dataa(Mux252),
	.datab(portB25),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~11_cout ),
	.combout(),
	.cout(\LessThan1~13_cout ));
// synopsys translate_off
defparam \LessThan1~13 .lut_mask = 16'h004D;
defparam \LessThan1~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N14
cycloneive_lcell_comb \LessThan1~15 (
// Equation(s):
// \LessThan1~15_cout  = CARRY((Mux242 & ((!\LessThan1~13_cout ) # (!\portB~51_combout ))) # (!Mux242 & (!\portB~51_combout  & !\LessThan1~13_cout )))

	.dataa(Mux242),
	.datab(portB24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~13_cout ),
	.combout(),
	.cout(\LessThan1~15_cout ));
// synopsys translate_off
defparam \LessThan1~15 .lut_mask = 16'h002B;
defparam \LessThan1~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N16
cycloneive_lcell_comb \LessThan1~17 (
// Equation(s):
// \LessThan1~17_cout  = CARRY((\portB~49_combout  & ((!\LessThan1~15_cout ) # (!Mux23))) # (!\portB~49_combout  & (!Mux23 & !\LessThan1~15_cout )))

	.dataa(portB23),
	.datab(Mux23),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~15_cout ),
	.combout(),
	.cout(\LessThan1~17_cout ));
// synopsys translate_off
defparam \LessThan1~17 .lut_mask = 16'h002B;
defparam \LessThan1~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N18
cycloneive_lcell_comb \LessThan1~19 (
// Equation(s):
// \LessThan1~19_cout  = CARRY((\portB~47_combout  & (Mux22 & !\LessThan1~17_cout )) # (!\portB~47_combout  & ((Mux22) # (!\LessThan1~17_cout ))))

	.dataa(portB22),
	.datab(Mux22),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~17_cout ),
	.combout(),
	.cout(\LessThan1~19_cout ));
// synopsys translate_off
defparam \LessThan1~19 .lut_mask = 16'h004D;
defparam \LessThan1~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N20
cycloneive_lcell_comb \LessThan1~21 (
// Equation(s):
// \LessThan1~21_cout  = CARRY((Mux21 & (\portB~45_combout  & !\LessThan1~19_cout )) # (!Mux21 & ((\portB~45_combout ) # (!\LessThan1~19_cout ))))

	.dataa(Mux21),
	.datab(portB21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~19_cout ),
	.combout(),
	.cout(\LessThan1~21_cout ));
// synopsys translate_off
defparam \LessThan1~21 .lut_mask = 16'h004D;
defparam \LessThan1~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N22
cycloneive_lcell_comb \LessThan1~23 (
// Equation(s):
// \LessThan1~23_cout  = CARRY((Mux20 & ((!\LessThan1~21_cout ) # (!\portB~43_combout ))) # (!Mux20 & (!\portB~43_combout  & !\LessThan1~21_cout )))

	.dataa(Mux20),
	.datab(portB20),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~21_cout ),
	.combout(),
	.cout(\LessThan1~23_cout ));
// synopsys translate_off
defparam \LessThan1~23 .lut_mask = 16'h002B;
defparam \LessThan1~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N24
cycloneive_lcell_comb \LessThan1~25 (
// Equation(s):
// \LessThan1~25_cout  = CARRY((\portB~41_combout  & ((!\LessThan1~23_cout ) # (!Mux19))) # (!\portB~41_combout  & (!Mux19 & !\LessThan1~23_cout )))

	.dataa(portB19),
	.datab(Mux19),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~23_cout ),
	.combout(),
	.cout(\LessThan1~25_cout ));
// synopsys translate_off
defparam \LessThan1~25 .lut_mask = 16'h002B;
defparam \LessThan1~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N26
cycloneive_lcell_comb \LessThan1~27 (
// Equation(s):
// \LessThan1~27_cout  = CARRY((\portB~39_combout  & (Mux18 & !\LessThan1~25_cout )) # (!\portB~39_combout  & ((Mux18) # (!\LessThan1~25_cout ))))

	.dataa(portB18),
	.datab(Mux18),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~25_cout ),
	.combout(),
	.cout(\LessThan1~27_cout ));
// synopsys translate_off
defparam \LessThan1~27 .lut_mask = 16'h004D;
defparam \LessThan1~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N28
cycloneive_lcell_comb \LessThan1~29 (
// Equation(s):
// \LessThan1~29_cout  = CARRY((Mux17 & (\portB~37_combout  & !\LessThan1~27_cout )) # (!Mux17 & ((\portB~37_combout ) # (!\LessThan1~27_cout ))))

	.dataa(Mux17),
	.datab(portB17),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~27_cout ),
	.combout(),
	.cout(\LessThan1~29_cout ));
// synopsys translate_off
defparam \LessThan1~29 .lut_mask = 16'h004D;
defparam \LessThan1~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N30
cycloneive_lcell_comb \LessThan1~31 (
// Equation(s):
// \LessThan1~31_cout  = CARRY((Mux16 & ((!\LessThan1~29_cout ) # (!\portB~35_combout ))) # (!Mux16 & (!\portB~35_combout  & !\LessThan1~29_cout )))

	.dataa(Mux16),
	.datab(portB16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~29_cout ),
	.combout(),
	.cout(\LessThan1~31_cout ));
// synopsys translate_off
defparam \LessThan1~31 .lut_mask = 16'h002B;
defparam \LessThan1~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N0
cycloneive_lcell_comb \LessThan1~33 (
// Equation(s):
// \LessThan1~33_cout  = CARRY((Mux15 & (\portB~33_combout  & !\LessThan1~31_cout )) # (!Mux15 & ((\portB~33_combout ) # (!\LessThan1~31_cout ))))

	.dataa(Mux15),
	.datab(portB15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~31_cout ),
	.combout(),
	.cout(\LessThan1~33_cout ));
// synopsys translate_off
defparam \LessThan1~33 .lut_mask = 16'h004D;
defparam \LessThan1~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N2
cycloneive_lcell_comb \LessThan1~35 (
// Equation(s):
// \LessThan1~35_cout  = CARRY((\portB~31_combout  & (Mux14 & !\LessThan1~33_cout )) # (!\portB~31_combout  & ((Mux14) # (!\LessThan1~33_cout ))))

	.dataa(portB14),
	.datab(Mux14),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~33_cout ),
	.combout(),
	.cout(\LessThan1~35_cout ));
// synopsys translate_off
defparam \LessThan1~35 .lut_mask = 16'h004D;
defparam \LessThan1~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N4
cycloneive_lcell_comb \LessThan1~37 (
// Equation(s):
// \LessThan1~37_cout  = CARRY((\portB~29_combout  & ((!\LessThan1~35_cout ) # (!Mux13))) # (!\portB~29_combout  & (!Mux13 & !\LessThan1~35_cout )))

	.dataa(portB13),
	.datab(Mux13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~35_cout ),
	.combout(),
	.cout(\LessThan1~37_cout ));
// synopsys translate_off
defparam \LessThan1~37 .lut_mask = 16'h002B;
defparam \LessThan1~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N6
cycloneive_lcell_comb \LessThan1~39 (
// Equation(s):
// \LessThan1~39_cout  = CARRY((Mux12 & ((!\LessThan1~37_cout ) # (!\portB~27_combout ))) # (!Mux12 & (!\portB~27_combout  & !\LessThan1~37_cout )))

	.dataa(Mux12),
	.datab(portB12),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~37_cout ),
	.combout(),
	.cout(\LessThan1~39_cout ));
// synopsys translate_off
defparam \LessThan1~39 .lut_mask = 16'h002B;
defparam \LessThan1~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N8
cycloneive_lcell_comb \LessThan1~41 (
// Equation(s):
// \LessThan1~41_cout  = CARRY((\portB~25_combout  & ((!\LessThan1~39_cout ) # (!Mux11))) # (!\portB~25_combout  & (!Mux11 & !\LessThan1~39_cout )))

	.dataa(portB11),
	.datab(Mux11),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~39_cout ),
	.combout(),
	.cout(\LessThan1~41_cout ));
// synopsys translate_off
defparam \LessThan1~41 .lut_mask = 16'h002B;
defparam \LessThan1~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N10
cycloneive_lcell_comb \LessThan1~43 (
// Equation(s):
// \LessThan1~43_cout  = CARRY((\portB~23_combout  & (Mux10 & !\LessThan1~41_cout )) # (!\portB~23_combout  & ((Mux10) # (!\LessThan1~41_cout ))))

	.dataa(portB10),
	.datab(Mux10),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~41_cout ),
	.combout(),
	.cout(\LessThan1~43_cout ));
// synopsys translate_off
defparam \LessThan1~43 .lut_mask = 16'h004D;
defparam \LessThan1~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N12
cycloneive_lcell_comb \LessThan1~45 (
// Equation(s):
// \LessThan1~45_cout  = CARRY((\portB~21_combout  & ((!\LessThan1~43_cout ) # (!Mux9))) # (!\portB~21_combout  & (!Mux9 & !\LessThan1~43_cout )))

	.dataa(portB9),
	.datab(Mux9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~43_cout ),
	.combout(),
	.cout(\LessThan1~45_cout ));
// synopsys translate_off
defparam \LessThan1~45 .lut_mask = 16'h002B;
defparam \LessThan1~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N14
cycloneive_lcell_comb \LessThan1~47 (
// Equation(s):
// \LessThan1~47_cout  = CARRY((Mux8 & ((!\LessThan1~45_cout ) # (!\portB~19_combout ))) # (!Mux8 & (!\portB~19_combout  & !\LessThan1~45_cout )))

	.dataa(Mux8),
	.datab(portB8),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~45_cout ),
	.combout(),
	.cout(\LessThan1~47_cout ));
// synopsys translate_off
defparam \LessThan1~47 .lut_mask = 16'h002B;
defparam \LessThan1~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N16
cycloneive_lcell_comb \LessThan1~49 (
// Equation(s):
// \LessThan1~49_cout  = CARRY((Mux72 & (\portB~17_combout  & !\LessThan1~47_cout )) # (!Mux72 & ((\portB~17_combout ) # (!\LessThan1~47_cout ))))

	.dataa(Mux72),
	.datab(portB7),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~47_cout ),
	.combout(),
	.cout(\LessThan1~49_cout ));
// synopsys translate_off
defparam \LessThan1~49 .lut_mask = 16'h004D;
defparam \LessThan1~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N18
cycloneive_lcell_comb \LessThan1~51 (
// Equation(s):
// \LessThan1~51_cout  = CARRY((\portB~15_combout  & (Mux6 & !\LessThan1~49_cout )) # (!\portB~15_combout  & ((Mux6) # (!\LessThan1~49_cout ))))

	.dataa(portB6),
	.datab(Mux6),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~49_cout ),
	.combout(),
	.cout(\LessThan1~51_cout ));
// synopsys translate_off
defparam \LessThan1~51 .lut_mask = 16'h004D;
defparam \LessThan1~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N20
cycloneive_lcell_comb \LessThan1~53 (
// Equation(s):
// \LessThan1~53_cout  = CARRY((Mux5 & (\portB~13_combout  & !\LessThan1~51_cout )) # (!Mux5 & ((\portB~13_combout ) # (!\LessThan1~51_cout ))))

	.dataa(Mux5),
	.datab(portB5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~51_cout ),
	.combout(),
	.cout(\LessThan1~53_cout ));
// synopsys translate_off
defparam \LessThan1~53 .lut_mask = 16'h004D;
defparam \LessThan1~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N22
cycloneive_lcell_comb \LessThan1~55 (
// Equation(s):
// \LessThan1~55_cout  = CARRY((\portB~11_combout  & (Mux4 & !\LessThan1~53_cout )) # (!\portB~11_combout  & ((Mux4) # (!\LessThan1~53_cout ))))

	.dataa(portB4),
	.datab(Mux4),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~53_cout ),
	.combout(),
	.cout(\LessThan1~55_cout ));
// synopsys translate_off
defparam \LessThan1~55 .lut_mask = 16'h004D;
defparam \LessThan1~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N24
cycloneive_lcell_comb \LessThan1~57 (
// Equation(s):
// \LessThan1~57_cout  = CARRY((Mux3 & (\portB~9_combout  & !\LessThan1~55_cout )) # (!Mux3 & ((\portB~9_combout ) # (!\LessThan1~55_cout ))))

	.dataa(Mux3),
	.datab(portB3),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~55_cout ),
	.combout(),
	.cout(\LessThan1~57_cout ));
// synopsys translate_off
defparam \LessThan1~57 .lut_mask = 16'h004D;
defparam \LessThan1~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N26
cycloneive_lcell_comb \LessThan1~59 (
// Equation(s):
// \LessThan1~59_cout  = CARRY((Mux2 & ((!\LessThan1~57_cout ) # (!\portB~7_combout ))) # (!Mux2 & (!\portB~7_combout  & !\LessThan1~57_cout )))

	.dataa(Mux2),
	.datab(portB2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~57_cout ),
	.combout(),
	.cout(\LessThan1~59_cout ));
// synopsys translate_off
defparam \LessThan1~59 .lut_mask = 16'h002B;
defparam \LessThan1~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N28
cycloneive_lcell_comb \LessThan1~61 (
// Equation(s):
// \LessThan1~61_cout  = CARRY((\portB~5_combout  & ((!\LessThan1~59_cout ) # (!Mux1))) # (!\portB~5_combout  & (!Mux1 & !\LessThan1~59_cout )))

	.dataa(portB1),
	.datab(Mux1),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~59_cout ),
	.combout(),
	.cout(\LessThan1~61_cout ));
// synopsys translate_off
defparam \LessThan1~61 .lut_mask = 16'h002B;
defparam \LessThan1~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N30
cycloneive_lcell_comb \LessThan1~62 (
// Equation(s):
// \LessThan1~62_combout  = (Mux0 & (\LessThan1~61_cout  & \portB~3_combout )) # (!Mux0 & ((\LessThan1~61_cout ) # (\portB~3_combout )))

	.dataa(gnd),
	.datab(Mux0),
	.datac(gnd),
	.datad(portB),
	.cin(\LessThan1~61_cout ),
	.combout(\LessThan1~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan1~62 .lut_mask = 16'hF330;
defparam \LessThan1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N8
cycloneive_lcell_comb \ShiftRight0~37 (
// Equation(s):
// \ShiftRight0~37_combout  = (!Mux302 & ((Mux312 & (\portB~63_combout )) # (!Mux312 & ((\portB~65_combout )))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB30),
	.datad(portB31),
	.cin(gnd),
	.combout(\ShiftRight0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~37 .lut_mask = 16'h3120;
defparam \ShiftRight0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N20
cycloneive_lcell_comb \ShiftRight0~38 (
// Equation(s):
// \ShiftRight0~38_combout  = (Mux312 & ((\portB~59_combout ))) # (!Mux312 & (\portB~61_combout ))

	.dataa(portB29),
	.datab(Mux312),
	.datac(gnd),
	.datad(portB28),
	.cin(gnd),
	.combout(\ShiftRight0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~38 .lut_mask = 16'hEE22;
defparam \ShiftRight0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N22
cycloneive_lcell_comb \ShiftRight0~39 (
// Equation(s):
// \ShiftRight0~39_combout  = (!Mux292 & ((\ShiftRight0~37_combout ) # ((Mux302 & \ShiftRight0~38_combout ))))

	.dataa(Mux292),
	.datab(Mux302),
	.datac(\ShiftRight0~37_combout ),
	.datad(\ShiftRight0~38_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~39 .lut_mask = 16'h5450;
defparam \ShiftRight0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N18
cycloneive_lcell_comb \ShiftRight0~40 (
// Equation(s):
// \ShiftRight0~40_combout  = (Mux302 & ((Mux312 & ((\portB~51_combout ))) # (!Mux312 & (\portB~53_combout ))))

	.dataa(portB25),
	.datab(Mux302),
	.datac(Mux312),
	.datad(portB24),
	.cin(gnd),
	.combout(\ShiftRight0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~40 .lut_mask = 16'hC808;
defparam \ShiftRight0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N24
cycloneive_lcell_comb \ShiftRight0~42 (
// Equation(s):
// \ShiftRight0~42_combout  = (\ShiftRight0~40_combout ) # ((\ShiftRight0~41_combout  & !Mux302))

	.dataa(\ShiftRight0~41_combout ),
	.datab(gnd),
	.datac(Mux302),
	.datad(\ShiftRight0~40_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~42 .lut_mask = 16'hFF0A;
defparam \ShiftRight0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N20
cycloneive_lcell_comb \ShiftRight0~43 (
// Equation(s):
// \ShiftRight0~43_combout  = (!Mux28 & ((\ShiftRight0~39_combout ) # ((Mux292 & \ShiftRight0~42_combout ))))

	.dataa(Mux28),
	.datab(Mux292),
	.datac(\ShiftRight0~39_combout ),
	.datad(\ShiftRight0~42_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~43 .lut_mask = 16'h5450;
defparam \ShiftRight0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N24
cycloneive_lcell_comb \ShiftRight0~123 (
// Equation(s):
// \ShiftRight0~123_combout  = (!Mux302 & ((dcifimemload_25 & ((!Mux31))) # (!dcifimemload_25 & (!Mux311))))

	.dataa(Mux311),
	.datab(Mux31),
	.datac(Mux302),
	.datad(dcifimemload_25),
	.cin(gnd),
	.combout(\ShiftRight0~123_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~123 .lut_mask = 16'h0305;
defparam \ShiftRight0~123 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N10
cycloneive_lcell_comb \ShiftRight0~44 (
// Equation(s):
// \ShiftRight0~44_combout  = (!Mux302 & (Mux312 & \portB~39_combout ))

	.dataa(gnd),
	.datab(Mux302),
	.datac(Mux312),
	.datad(portB18),
	.cin(gnd),
	.combout(\ShiftRight0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~44 .lut_mask = 16'h3000;
defparam \ShiftRight0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N18
cycloneive_lcell_comb \ShiftRight0~45 (
// Equation(s):
// \ShiftRight0~45_combout  = (Mux302 & ((Mux312 & ((\portB~35_combout ))) # (!Mux312 & (\portB~37_combout ))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB17),
	.datad(portB16),
	.cin(gnd),
	.combout(\ShiftRight0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~45 .lut_mask = 16'hC840;
defparam \ShiftRight0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N0
cycloneive_lcell_comb \ShiftRight0~46 (
// Equation(s):
// \ShiftRight0~46_combout  = (\ShiftRight0~44_combout ) # ((\ShiftRight0~45_combout ) # ((\portB~41_combout  & \ShiftRight0~123_combout )))

	.dataa(portB19),
	.datab(\ShiftRight0~123_combout ),
	.datac(\ShiftRight0~44_combout ),
	.datad(\ShiftRight0~45_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~46 .lut_mask = 16'hFFF8;
defparam \ShiftRight0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N18
cycloneive_lcell_comb \ShiftRight0~47 (
// Equation(s):
// \ShiftRight0~47_combout  = (Mux302 & ((Mux312 & ((\portB~43_combout ))) # (!Mux312 & (\portB~45_combout )))) # (!Mux302 & (((Mux312))))

	.dataa(portB21),
	.datab(portB20),
	.datac(Mux302),
	.datad(Mux312),
	.cin(gnd),
	.combout(\ShiftRight0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~47 .lut_mask = 16'hCFA0;
defparam \ShiftRight0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N24
cycloneive_lcell_comb \ShiftRight0~48 (
// Equation(s):
// \ShiftRight0~48_combout  = (Mux302 & (((\ShiftRight0~47_combout )))) # (!Mux302 & ((\ShiftRight0~47_combout  & ((\portB~47_combout ))) # (!\ShiftRight0~47_combout  & (\portB~49_combout ))))

	.dataa(portB23),
	.datab(Mux302),
	.datac(portB22),
	.datad(\ShiftRight0~47_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~48 .lut_mask = 16'hFC22;
defparam \ShiftRight0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N30
cycloneive_lcell_comb \ShiftRight0~49 (
// Equation(s):
// \ShiftRight0~49_combout  = (Mux28 & ((Mux292 & (\ShiftRight0~46_combout )) # (!Mux292 & ((\ShiftRight0~48_combout )))))

	.dataa(Mux28),
	.datab(\ShiftRight0~46_combout ),
	.datac(\ShiftRight0~48_combout ),
	.datad(Mux292),
	.cin(gnd),
	.combout(\ShiftRight0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~49 .lut_mask = 16'h88A0;
defparam \ShiftRight0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N16
cycloneive_lcell_comb \ShiftRight0~35 (
// Equation(s):
// \ShiftRight0~35_combout  = (Mux302 & ((Mux312 & (\portB~27_combout )) # (!Mux312 & ((\portB~29_combout )))))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB12),
	.datad(portB13),
	.cin(gnd),
	.combout(\ShiftRight0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~35 .lut_mask = 16'hA280;
defparam \ShiftRight0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N28
cycloneive_lcell_comb \ShiftRight0~31 (
// Equation(s):
// \ShiftRight0~31_combout  = (!Mux302 & (\portB~23_combout  & Mux312))

	.dataa(gnd),
	.datab(Mux302),
	.datac(portB10),
	.datad(Mux312),
	.cin(gnd),
	.combout(\ShiftRight0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~31 .lut_mask = 16'h3000;
defparam \ShiftRight0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N22
cycloneive_lcell_comb \ShiftRight0~32 (
// Equation(s):
// \ShiftRight0~32_combout  = (Mux302 & ((Mux312 & ((\portB~19_combout ))) # (!Mux312 & (\portB~21_combout ))))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB9),
	.datad(portB8),
	.cin(gnd),
	.combout(\ShiftRight0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~32 .lut_mask = 16'hA820;
defparam \ShiftRight0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N12
cycloneive_lcell_comb \ShiftRight0~33 (
// Equation(s):
// \ShiftRight0~33_combout  = (\ShiftRight0~31_combout ) # ((\ShiftRight0~32_combout ) # ((\portB~25_combout  & \ShiftRight0~123_combout )))

	.dataa(portB11),
	.datab(\ShiftRight0~31_combout ),
	.datac(\ShiftRight0~32_combout ),
	.datad(\ShiftRight0~123_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~33 .lut_mask = 16'hFEFC;
defparam \ShiftRight0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N6
cycloneive_lcell_comb \Selector23~2 (
// Equation(s):
// \Selector23~2_combout  = (Mux292 & (((\ShiftRight0~33_combout )))) # (!Mux292 & ((\ShiftRight0~34_combout ) # ((\ShiftRight0~35_combout ))))

	.dataa(\ShiftRight0~34_combout ),
	.datab(\ShiftRight0~35_combout ),
	.datac(Mux292),
	.datad(\ShiftRight0~33_combout ),
	.cin(gnd),
	.combout(\Selector23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~2 .lut_mask = 16'hFE0E;
defparam \Selector23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N4
cycloneive_lcell_comb \ShiftRight0~24 (
// Equation(s):
// \ShiftRight0~24_combout  = (!Mux302 & ((Mux312 & ((\portB~7_combout ))) # (!Mux312 & (\portB~9_combout ))))

	.dataa(portB3),
	.datab(Mux312),
	.datac(Mux302),
	.datad(portB2),
	.cin(gnd),
	.combout(\ShiftRight0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~24 .lut_mask = 16'h0E02;
defparam \ShiftRight0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N10
cycloneive_lcell_comb \ShiftRight0~25 (
// Equation(s):
// \ShiftRight0~25_combout  = (Mux312 & (\portB~3_combout )) # (!Mux312 & ((\portB~5_combout )))

	.dataa(gnd),
	.datab(Mux312),
	.datac(portB),
	.datad(portB1),
	.cin(gnd),
	.combout(\ShiftRight0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~25 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N24
cycloneive_lcell_comb \ShiftRight0~26 (
// Equation(s):
// \ShiftRight0~26_combout  = (\ShiftRight0~24_combout ) # ((Mux302 & \ShiftRight0~25_combout ))

	.dataa(gnd),
	.datab(Mux302),
	.datac(\ShiftRight0~24_combout ),
	.datad(\ShiftRight0~25_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~26 .lut_mask = 16'hFCF0;
defparam \ShiftRight0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N24
cycloneive_lcell_comb \ShiftRight0~122 (
// Equation(s):
// \ShiftRight0~122_combout  = (!Mux312 & ((dcifimemload_25 & ((Mux30))) # (!dcifimemload_25 & (Mux301))))

	.dataa(dcifimemload_25),
	.datab(Mux301),
	.datac(Mux312),
	.datad(Mux30),
	.cin(gnd),
	.combout(\ShiftRight0~122_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~122 .lut_mask = 16'h0E04;
defparam \ShiftRight0~122 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N20
cycloneive_lcell_comb \ShiftRight0~27 (
// Equation(s):
// \ShiftRight0~27_combout  = (Mux312 & (Mux302 & (\portB~11_combout ))) # (!Mux312 & (!Mux302 & ((\portB~17_combout ))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB4),
	.datad(portB7),
	.cin(gnd),
	.combout(\ShiftRight0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~27 .lut_mask = 16'h9180;
defparam \ShiftRight0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N10
cycloneive_lcell_comb \ShiftRight0~28 (
// Equation(s):
// \ShiftRight0~28_combout  = (\ShiftRight0~27_combout ) # ((Mux312 & (!Mux302 & \portB~15_combout )))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB6),
	.datad(\ShiftRight0~27_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~28 .lut_mask = 16'hFF20;
defparam \ShiftRight0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N24
cycloneive_lcell_comb \ShiftRight0~29 (
// Equation(s):
// \ShiftRight0~29_combout  = (\ShiftRight0~28_combout ) # ((\ShiftRight0~122_combout  & \portB~13_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~122_combout ),
	.datac(portB5),
	.datad(\ShiftRight0~28_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~29 .lut_mask = 16'hFFC0;
defparam \ShiftRight0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N6
cycloneive_lcell_comb \ShiftRight0~30 (
// Equation(s):
// \ShiftRight0~30_combout  = (Mux292 & (\ShiftRight0~26_combout )) # (!Mux292 & ((\ShiftRight0~29_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~26_combout ),
	.datac(Mux292),
	.datad(\ShiftRight0~29_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~30 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N0
cycloneive_lcell_comb \ShiftRight0~36 (
// Equation(s):
// \ShiftRight0~36_combout  = (Mux28 & ((\ShiftRight0~30_combout ))) # (!Mux28 & (\Selector23~2_combout ))

	.dataa(\Selector23~2_combout ),
	.datab(gnd),
	.datac(Mux28),
	.datad(\ShiftRight0~30_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~36 .lut_mask = 16'hFA0A;
defparam \ShiftRight0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N18
cycloneive_lcell_comb \Selector0~13 (
// Equation(s):
// \Selector0~13_combout  = (cuifALUOP_0 & (!cuifALUOP_3 & (!cuifALUOP_1 & !cuifALUOP_2)))

	.dataa(cuifALUOP_0),
	.datab(cuifALUOP_3),
	.datac(cuifALUOP_1),
	.datad(cuifALUOP_2),
	.cin(gnd),
	.combout(\Selector0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~13 .lut_mask = 16'h0002;
defparam \Selector0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N20
cycloneive_lcell_comb \Selector0~20 (
// Equation(s):
// \Selector0~20_combout  = (cuifALUOP_0 & (!cuifALUOP_1 & (!cuifALUOP_3 & !cuifALUOP_2)))

	.dataa(cuifALUOP_0),
	.datab(cuifALUOP_1),
	.datac(cuifALUOP_3),
	.datad(cuifALUOP_2),
	.cin(gnd),
	.combout(\Selector0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~20 .lut_mask = 16'h0002;
defparam \Selector0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N2
cycloneive_lcell_comb \Selector0~14 (
// Equation(s):
// \Selector0~14_combout  = (cuifALUOP_0 & (cuifALUOP_1 & (!cuifALUOP_3 & !cuifALUOP_2)))

	.dataa(cuifALUOP_0),
	.datab(cuifALUOP_1),
	.datac(cuifALUOP_3),
	.datad(cuifALUOP_2),
	.cin(gnd),
	.combout(\Selector0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~14 .lut_mask = 16'h0008;
defparam \Selector0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N2
cycloneive_lcell_comb \Add1~2 (
// Equation(s):
// \Add1~2_combout  = (\portB~63_combout  & ((Mux302 & (!\Add1~1 )) # (!Mux302 & ((\Add1~1 ) # (GND))))) # (!\portB~63_combout  & ((Mux302 & (\Add1~1  & VCC)) # (!Mux302 & (!\Add1~1 ))))
// \Add1~3  = CARRY((\portB~63_combout  & ((!\Add1~1 ) # (!Mux302))) # (!\portB~63_combout  & (!Mux302 & !\Add1~1 )))

	.dataa(portB30),
	.datab(Mux302),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h692B;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N4
cycloneive_lcell_comb \Add1~4 (
// Equation(s):
// \Add1~4_combout  = ((Mux292 $ (\portB~61_combout  $ (\Add1~3 )))) # (GND)
// \Add1~5  = CARRY((Mux292 & ((!\Add1~3 ) # (!\portB~61_combout ))) # (!Mux292 & (!\portB~61_combout  & !\Add1~3 )))

	.dataa(Mux292),
	.datab(portB29),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'h962B;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N6
cycloneive_lcell_comb \Add1~6 (
// Equation(s):
// \Add1~6_combout  = (Mux28 & ((\portB~59_combout  & (!\Add1~5 )) # (!\portB~59_combout  & (\Add1~5  & VCC)))) # (!Mux28 & ((\portB~59_combout  & ((\Add1~5 ) # (GND))) # (!\portB~59_combout  & (!\Add1~5 ))))
// \Add1~7  = CARRY((Mux28 & (\portB~59_combout  & !\Add1~5 )) # (!Mux28 & ((\portB~59_combout ) # (!\Add1~5 ))))

	.dataa(Mux28),
	.datab(portB28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h694D;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N8
cycloneive_lcell_comb \Add1~8 (
// Equation(s):
// \Add1~8_combout  = ((\portB~57_combout  $ (Mux272 $ (\Add1~7 )))) # (GND)
// \Add1~9  = CARRY((\portB~57_combout  & (Mux272 & !\Add1~7 )) # (!\portB~57_combout  & ((Mux272) # (!\Add1~7 ))))

	.dataa(portB27),
	.datab(Mux272),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'h964D;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N10
cycloneive_lcell_comb \Add1~10 (
// Equation(s):
// \Add1~10_combout  = (Mux26 & ((\portB~55_combout  & (!\Add1~9 )) # (!\portB~55_combout  & (\Add1~9  & VCC)))) # (!Mux26 & ((\portB~55_combout  & ((\Add1~9 ) # (GND))) # (!\portB~55_combout  & (!\Add1~9 ))))
// \Add1~11  = CARRY((Mux26 & (\portB~55_combout  & !\Add1~9 )) # (!Mux26 & ((\portB~55_combout ) # (!\Add1~9 ))))

	.dataa(Mux26),
	.datab(portB26),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h694D;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N12
cycloneive_lcell_comb \Add1~12 (
// Equation(s):
// \Add1~12_combout  = ((\portB~53_combout  $ (Mux252 $ (\Add1~11 )))) # (GND)
// \Add1~13  = CARRY((\portB~53_combout  & (Mux252 & !\Add1~11 )) # (!\portB~53_combout  & ((Mux252) # (!\Add1~11 ))))

	.dataa(portB25),
	.datab(Mux252),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
// synopsys translate_off
defparam \Add1~12 .lut_mask = 16'h964D;
defparam \Add1~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N14
cycloneive_lcell_comb \Add1~14 (
// Equation(s):
// \Add1~14_combout  = (\portB~51_combout  & ((Mux242 & (!\Add1~13 )) # (!Mux242 & ((\Add1~13 ) # (GND))))) # (!\portB~51_combout  & ((Mux242 & (\Add1~13  & VCC)) # (!Mux242 & (!\Add1~13 ))))
// \Add1~15  = CARRY((\portB~51_combout  & ((!\Add1~13 ) # (!Mux242))) # (!\portB~51_combout  & (!Mux242 & !\Add1~13 )))

	.dataa(portB24),
	.datab(Mux242),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
// synopsys translate_off
defparam \Add1~14 .lut_mask = 16'h692B;
defparam \Add1~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N16
cycloneive_lcell_comb \Add1~16 (
// Equation(s):
// \Add1~16_combout  = ((Mux23 $ (\portB~49_combout  $ (\Add1~15 )))) # (GND)
// \Add1~17  = CARRY((Mux23 & ((!\Add1~15 ) # (!\portB~49_combout ))) # (!Mux23 & (!\portB~49_combout  & !\Add1~15 )))

	.dataa(Mux23),
	.datab(portB23),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout(\Add1~17 ));
// synopsys translate_off
defparam \Add1~16 .lut_mask = 16'h962B;
defparam \Add1~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N18
cycloneive_lcell_comb \Add1~18 (
// Equation(s):
// \Add1~18_combout  = (Mux22 & ((\portB~47_combout  & (!\Add1~17 )) # (!\portB~47_combout  & (\Add1~17  & VCC)))) # (!Mux22 & ((\portB~47_combout  & ((\Add1~17 ) # (GND))) # (!\portB~47_combout  & (!\Add1~17 ))))
// \Add1~19  = CARRY((Mux22 & (\portB~47_combout  & !\Add1~17 )) # (!Mux22 & ((\portB~47_combout ) # (!\Add1~17 ))))

	.dataa(Mux22),
	.datab(portB22),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~17 ),
	.combout(\Add1~18_combout ),
	.cout(\Add1~19 ));
// synopsys translate_off
defparam \Add1~18 .lut_mask = 16'h694D;
defparam \Add1~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N20
cycloneive_lcell_comb \Add1~20 (
// Equation(s):
// \Add1~20_combout  = ((\portB~45_combout  $ (Mux21 $ (\Add1~19 )))) # (GND)
// \Add1~21  = CARRY((\portB~45_combout  & (Mux21 & !\Add1~19 )) # (!\portB~45_combout  & ((Mux21) # (!\Add1~19 ))))

	.dataa(portB21),
	.datab(Mux21),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~19 ),
	.combout(\Add1~20_combout ),
	.cout(\Add1~21 ));
// synopsys translate_off
defparam \Add1~20 .lut_mask = 16'h964D;
defparam \Add1~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N22
cycloneive_lcell_comb \Add1~22 (
// Equation(s):
// \Add1~22_combout  = (\portB~43_combout  & ((Mux20 & (!\Add1~21 )) # (!Mux20 & ((\Add1~21 ) # (GND))))) # (!\portB~43_combout  & ((Mux20 & (\Add1~21  & VCC)) # (!Mux20 & (!\Add1~21 ))))
// \Add1~23  = CARRY((\portB~43_combout  & ((!\Add1~21 ) # (!Mux20))) # (!\portB~43_combout  & (!Mux20 & !\Add1~21 )))

	.dataa(portB20),
	.datab(Mux20),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~21 ),
	.combout(\Add1~22_combout ),
	.cout(\Add1~23 ));
// synopsys translate_off
defparam \Add1~22 .lut_mask = 16'h692B;
defparam \Add1~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N24
cycloneive_lcell_comb \Add1~24 (
// Equation(s):
// \Add1~24_combout  = ((Mux19 $ (\portB~41_combout  $ (\Add1~23 )))) # (GND)
// \Add1~25  = CARRY((Mux19 & ((!\Add1~23 ) # (!\portB~41_combout ))) # (!Mux19 & (!\portB~41_combout  & !\Add1~23 )))

	.dataa(Mux19),
	.datab(portB19),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~23 ),
	.combout(\Add1~24_combout ),
	.cout(\Add1~25 ));
// synopsys translate_off
defparam \Add1~24 .lut_mask = 16'h962B;
defparam \Add1~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N28
cycloneive_lcell_comb \Add1~28 (
// Equation(s):
// \Add1~28_combout  = ((Mux17 $ (\portB~37_combout  $ (\Add1~27 )))) # (GND)
// \Add1~29  = CARRY((Mux17 & ((!\Add1~27 ) # (!\portB~37_combout ))) # (!Mux17 & (!\portB~37_combout  & !\Add1~27 )))

	.dataa(Mux17),
	.datab(portB17),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~27 ),
	.combout(\Add1~28_combout ),
	.cout(\Add1~29 ));
// synopsys translate_off
defparam \Add1~28 .lut_mask = 16'h962B;
defparam \Add1~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N30
cycloneive_lcell_comb \Add1~30 (
// Equation(s):
// \Add1~30_combout  = (\portB~35_combout  & ((Mux16 & (!\Add1~29 )) # (!Mux16 & ((\Add1~29 ) # (GND))))) # (!\portB~35_combout  & ((Mux16 & (\Add1~29  & VCC)) # (!Mux16 & (!\Add1~29 ))))
// \Add1~31  = CARRY((\portB~35_combout  & ((!\Add1~29 ) # (!Mux16))) # (!\portB~35_combout  & (!Mux16 & !\Add1~29 )))

	.dataa(portB16),
	.datab(Mux16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~29 ),
	.combout(\Add1~30_combout ),
	.cout(\Add1~31 ));
// synopsys translate_off
defparam \Add1~30 .lut_mask = 16'h692B;
defparam \Add1~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N0
cycloneive_lcell_comb \Add1~32 (
// Equation(s):
// \Add1~32_combout  = ((\portB~33_combout  $ (Mux15 $ (\Add1~31 )))) # (GND)
// \Add1~33  = CARRY((\portB~33_combout  & (Mux15 & !\Add1~31 )) # (!\portB~33_combout  & ((Mux15) # (!\Add1~31 ))))

	.dataa(portB15),
	.datab(Mux15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~31 ),
	.combout(\Add1~32_combout ),
	.cout(\Add1~33 ));
// synopsys translate_off
defparam \Add1~32 .lut_mask = 16'h964D;
defparam \Add1~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N2
cycloneive_lcell_comb \Add1~34 (
// Equation(s):
// \Add1~34_combout  = (\portB~31_combout  & ((Mux14 & (!\Add1~33 )) # (!Mux14 & ((\Add1~33 ) # (GND))))) # (!\portB~31_combout  & ((Mux14 & (\Add1~33  & VCC)) # (!Mux14 & (!\Add1~33 ))))
// \Add1~35  = CARRY((\portB~31_combout  & ((!\Add1~33 ) # (!Mux14))) # (!\portB~31_combout  & (!Mux14 & !\Add1~33 )))

	.dataa(portB14),
	.datab(Mux14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~33 ),
	.combout(\Add1~34_combout ),
	.cout(\Add1~35 ));
// synopsys translate_off
defparam \Add1~34 .lut_mask = 16'h692B;
defparam \Add1~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N4
cycloneive_lcell_comb \Add1~36 (
// Equation(s):
// \Add1~36_combout  = ((\portB~29_combout  $ (Mux13 $ (\Add1~35 )))) # (GND)
// \Add1~37  = CARRY((\portB~29_combout  & (Mux13 & !\Add1~35 )) # (!\portB~29_combout  & ((Mux13) # (!\Add1~35 ))))

	.dataa(portB13),
	.datab(Mux13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~35 ),
	.combout(\Add1~36_combout ),
	.cout(\Add1~37 ));
// synopsys translate_off
defparam \Add1~36 .lut_mask = 16'h964D;
defparam \Add1~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N6
cycloneive_lcell_comb \Add1~38 (
// Equation(s):
// \Add1~38_combout  = (\portB~27_combout  & ((Mux12 & (!\Add1~37 )) # (!Mux12 & ((\Add1~37 ) # (GND))))) # (!\portB~27_combout  & ((Mux12 & (\Add1~37  & VCC)) # (!Mux12 & (!\Add1~37 ))))
// \Add1~39  = CARRY((\portB~27_combout  & ((!\Add1~37 ) # (!Mux12))) # (!\portB~27_combout  & (!Mux12 & !\Add1~37 )))

	.dataa(portB12),
	.datab(Mux12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~37 ),
	.combout(\Add1~38_combout ),
	.cout(\Add1~39 ));
// synopsys translate_off
defparam \Add1~38 .lut_mask = 16'h692B;
defparam \Add1~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N8
cycloneive_lcell_comb \Add1~40 (
// Equation(s):
// \Add1~40_combout  = ((Mux11 $ (\portB~25_combout  $ (\Add1~39 )))) # (GND)
// \Add1~41  = CARRY((Mux11 & ((!\Add1~39 ) # (!\portB~25_combout ))) # (!Mux11 & (!\portB~25_combout  & !\Add1~39 )))

	.dataa(Mux11),
	.datab(portB11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~39 ),
	.combout(\Add1~40_combout ),
	.cout(\Add1~41 ));
// synopsys translate_off
defparam \Add1~40 .lut_mask = 16'h962B;
defparam \Add1~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N10
cycloneive_lcell_comb \Add1~42 (
// Equation(s):
// \Add1~42_combout  = (\portB~23_combout  & ((Mux10 & (!\Add1~41 )) # (!Mux10 & ((\Add1~41 ) # (GND))))) # (!\portB~23_combout  & ((Mux10 & (\Add1~41  & VCC)) # (!Mux10 & (!\Add1~41 ))))
// \Add1~43  = CARRY((\portB~23_combout  & ((!\Add1~41 ) # (!Mux10))) # (!\portB~23_combout  & (!Mux10 & !\Add1~41 )))

	.dataa(portB10),
	.datab(Mux10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~41 ),
	.combout(\Add1~42_combout ),
	.cout(\Add1~43 ));
// synopsys translate_off
defparam \Add1~42 .lut_mask = 16'h692B;
defparam \Add1~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N12
cycloneive_lcell_comb \Add1~44 (
// Equation(s):
// \Add1~44_combout  = ((\portB~21_combout  $ (Mux9 $ (\Add1~43 )))) # (GND)
// \Add1~45  = CARRY((\portB~21_combout  & (Mux9 & !\Add1~43 )) # (!\portB~21_combout  & ((Mux9) # (!\Add1~43 ))))

	.dataa(portB9),
	.datab(Mux9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~43 ),
	.combout(\Add1~44_combout ),
	.cout(\Add1~45 ));
// synopsys translate_off
defparam \Add1~44 .lut_mask = 16'h964D;
defparam \Add1~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N14
cycloneive_lcell_comb \Add1~46 (
// Equation(s):
// \Add1~46_combout  = (Mux8 & ((\portB~19_combout  & (!\Add1~45 )) # (!\portB~19_combout  & (\Add1~45  & VCC)))) # (!Mux8 & ((\portB~19_combout  & ((\Add1~45 ) # (GND))) # (!\portB~19_combout  & (!\Add1~45 ))))
// \Add1~47  = CARRY((Mux8 & (\portB~19_combout  & !\Add1~45 )) # (!Mux8 & ((\portB~19_combout ) # (!\Add1~45 ))))

	.dataa(Mux8),
	.datab(portB8),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~45 ),
	.combout(\Add1~46_combout ),
	.cout(\Add1~47 ));
// synopsys translate_off
defparam \Add1~46 .lut_mask = 16'h694D;
defparam \Add1~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N16
cycloneive_lcell_comb \Add1~48 (
// Equation(s):
// \Add1~48_combout  = ((Mux72 $ (\portB~17_combout  $ (\Add1~47 )))) # (GND)
// \Add1~49  = CARRY((Mux72 & ((!\Add1~47 ) # (!\portB~17_combout ))) # (!Mux72 & (!\portB~17_combout  & !\Add1~47 )))

	.dataa(Mux72),
	.datab(portB7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~47 ),
	.combout(\Add1~48_combout ),
	.cout(\Add1~49 ));
// synopsys translate_off
defparam \Add1~48 .lut_mask = 16'h962B;
defparam \Add1~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N18
cycloneive_lcell_comb \Add1~50 (
// Equation(s):
// \Add1~50_combout  = (\portB~15_combout  & ((Mux6 & (!\Add1~49 )) # (!Mux6 & ((\Add1~49 ) # (GND))))) # (!\portB~15_combout  & ((Mux6 & (\Add1~49  & VCC)) # (!Mux6 & (!\Add1~49 ))))
// \Add1~51  = CARRY((\portB~15_combout  & ((!\Add1~49 ) # (!Mux6))) # (!\portB~15_combout  & (!Mux6 & !\Add1~49 )))

	.dataa(portB6),
	.datab(Mux6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~49 ),
	.combout(\Add1~50_combout ),
	.cout(\Add1~51 ));
// synopsys translate_off
defparam \Add1~50 .lut_mask = 16'h692B;
defparam \Add1~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N20
cycloneive_lcell_comb \Add1~52 (
// Equation(s):
// \Add1~52_combout  = ((Mux5 $ (\portB~13_combout  $ (\Add1~51 )))) # (GND)
// \Add1~53  = CARRY((Mux5 & ((!\Add1~51 ) # (!\portB~13_combout ))) # (!Mux5 & (!\portB~13_combout  & !\Add1~51 )))

	.dataa(Mux5),
	.datab(portB5),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~51 ),
	.combout(\Add1~52_combout ),
	.cout(\Add1~53 ));
// synopsys translate_off
defparam \Add1~52 .lut_mask = 16'h962B;
defparam \Add1~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N22
cycloneive_lcell_comb \Add1~54 (
// Equation(s):
// \Add1~54_combout  = (Mux4 & ((\portB~11_combout  & (!\Add1~53 )) # (!\portB~11_combout  & (\Add1~53  & VCC)))) # (!Mux4 & ((\portB~11_combout  & ((\Add1~53 ) # (GND))) # (!\portB~11_combout  & (!\Add1~53 ))))
// \Add1~55  = CARRY((Mux4 & (\portB~11_combout  & !\Add1~53 )) # (!Mux4 & ((\portB~11_combout ) # (!\Add1~53 ))))

	.dataa(Mux4),
	.datab(portB4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~53 ),
	.combout(\Add1~54_combout ),
	.cout(\Add1~55 ));
// synopsys translate_off
defparam \Add1~54 .lut_mask = 16'h694D;
defparam \Add1~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N24
cycloneive_lcell_comb \Add1~56 (
// Equation(s):
// \Add1~56_combout  = ((\portB~9_combout  $ (Mux3 $ (\Add1~55 )))) # (GND)
// \Add1~57  = CARRY((\portB~9_combout  & (Mux3 & !\Add1~55 )) # (!\portB~9_combout  & ((Mux3) # (!\Add1~55 ))))

	.dataa(portB3),
	.datab(Mux3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~55 ),
	.combout(\Add1~56_combout ),
	.cout(\Add1~57 ));
// synopsys translate_off
defparam \Add1~56 .lut_mask = 16'h964D;
defparam \Add1~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N26
cycloneive_lcell_comb \Add1~58 (
// Equation(s):
// \Add1~58_combout  = (Mux2 & ((\portB~7_combout  & (!\Add1~57 )) # (!\portB~7_combout  & (\Add1~57  & VCC)))) # (!Mux2 & ((\portB~7_combout  & ((\Add1~57 ) # (GND))) # (!\portB~7_combout  & (!\Add1~57 ))))
// \Add1~59  = CARRY((Mux2 & (\portB~7_combout  & !\Add1~57 )) # (!Mux2 & ((\portB~7_combout ) # (!\Add1~57 ))))

	.dataa(Mux2),
	.datab(portB2),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~57 ),
	.combout(\Add1~58_combout ),
	.cout(\Add1~59 ));
// synopsys translate_off
defparam \Add1~58 .lut_mask = 16'h694D;
defparam \Add1~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N28
cycloneive_lcell_comb \Add1~60 (
// Equation(s):
// \Add1~60_combout  = ((Mux1 $ (\portB~5_combout  $ (\Add1~59 )))) # (GND)
// \Add1~61  = CARRY((Mux1 & ((!\Add1~59 ) # (!\portB~5_combout ))) # (!Mux1 & (!\portB~5_combout  & !\Add1~59 )))

	.dataa(Mux1),
	.datab(portB1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~59 ),
	.combout(\Add1~60_combout ),
	.cout(\Add1~61 ));
// synopsys translate_off
defparam \Add1~60 .lut_mask = 16'h962B;
defparam \Add1~60 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N30
cycloneive_lcell_comb \Add1~62 (
// Equation(s):
// \Add1~62_combout  = Mux0 $ (\Add1~61  $ (!\portB~3_combout ))

	.dataa(Mux0),
	.datab(gnd),
	.datac(gnd),
	.datad(portB),
	.cin(\Add1~61 ),
	.combout(\Add1~62_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~62 .lut_mask = 16'h5AA5;
defparam \Add1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N26
cycloneive_lcell_comb \Selector0~17 (
// Equation(s):
// \Selector0~17_combout  = (cuifALUOP_2 & (cuifALUOP_0 & (!cuifALUOP_3 & !cuifALUOP_1)))

	.dataa(cuifALUOP_2),
	.datab(cuifALUOP_0),
	.datac(cuifALUOP_3),
	.datad(cuifALUOP_1),
	.cin(gnd),
	.combout(\Selector0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~17 .lut_mask = 16'h0008;
defparam \Selector0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N30
cycloneive_lcell_comb \Selector0~28 (
// Equation(s):
// \Selector0~28_combout  = (Mux0 & (((\Selector0~17_combout )))) # (!Mux0 & (\Selector0~27_combout  & ((!\portB~3_combout ))))

	.dataa(\Selector0~27_combout ),
	.datab(\Selector0~17_combout ),
	.datac(portB),
	.datad(Mux0),
	.cin(gnd),
	.combout(\Selector0~28_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~28 .lut_mask = 16'hCC0A;
defparam \Selector0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N28
cycloneive_lcell_comb \Selector0~15 (
// Equation(s):
// \Selector0~15_combout  = (cuifALUOP_2 & (cuifALUOP_1 & (!cuifALUOP_3 & !cuifALUOP_0)))

	.dataa(cuifALUOP_2),
	.datab(cuifALUOP_1),
	.datac(cuifALUOP_3),
	.datad(cuifALUOP_0),
	.cin(gnd),
	.combout(\Selector0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~15 .lut_mask = 16'h0008;
defparam \Selector0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N26
cycloneive_lcell_comb \Selector0~16 (
// Equation(s):
// \Selector0~16_combout  = (\Selector0~15_combout  & (\portB~3_combout  $ (Mux0)))

	.dataa(gnd),
	.datab(\Selector0~15_combout ),
	.datac(portB),
	.datad(Mux0),
	.cin(gnd),
	.combout(\Selector0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~16 .lut_mask = 16'h0CC0;
defparam \Selector0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N22
cycloneive_lcell_comb \ShiftLeft0~12 (
// Equation(s):
// \ShiftLeft0~12_combout  = (\portB~23_combout  & ((\ShiftRight0~122_combout ) # ((\ShiftRight0~123_combout  & \portB~19_combout )))) # (!\portB~23_combout  & (\ShiftRight0~123_combout  & ((\portB~19_combout ))))

	.dataa(portB10),
	.datab(\ShiftRight0~123_combout ),
	.datac(\ShiftRight0~122_combout ),
	.datad(portB8),
	.cin(gnd),
	.combout(\ShiftLeft0~12_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~12 .lut_mask = 16'hECA0;
defparam \ShiftLeft0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N28
cycloneive_lcell_comb \ShiftLeft0~11 (
// Equation(s):
// \ShiftLeft0~11_combout  = (Mux312 & ((Mux302 & (\portB~25_combout )) # (!Mux302 & ((\portB~21_combout )))))

	.dataa(Mux302),
	.datab(portB11),
	.datac(Mux312),
	.datad(portB9),
	.cin(gnd),
	.combout(\ShiftLeft0~11_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~11 .lut_mask = 16'hD080;
defparam \ShiftLeft0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N4
cycloneive_lcell_comb \ShiftLeft0~13 (
// Equation(s):
// \ShiftLeft0~13_combout  = (\ShiftLeft0~12_combout ) # (\ShiftLeft0~11_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftLeft0~12_combout ),
	.datad(\ShiftLeft0~11_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~13_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~13 .lut_mask = 16'hFFF0;
defparam \ShiftLeft0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N0
cycloneive_lcell_comb \ShiftLeft0~8 (
// Equation(s):
// \ShiftLeft0~8_combout  = (Mux312 & ((Mux302 & (\portB~33_combout )) # (!Mux302 & ((\portB~29_combout )))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB15),
	.datad(portB13),
	.cin(gnd),
	.combout(\ShiftLeft0~8_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~8 .lut_mask = 16'hA280;
defparam \ShiftLeft0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N2
cycloneive_lcell_comb \ShiftLeft0~9 (
// Equation(s):
// \ShiftLeft0~9_combout  = (\portB~27_combout  & ((\ShiftRight0~123_combout ) # ((\portB~31_combout  & \ShiftRight0~122_combout )))) # (!\portB~27_combout  & (\portB~31_combout  & (\ShiftRight0~122_combout )))

	.dataa(portB12),
	.datab(portB14),
	.datac(\ShiftRight0~122_combout ),
	.datad(\ShiftRight0~123_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~9_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~9 .lut_mask = 16'hEAC0;
defparam \ShiftLeft0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N2
cycloneive_lcell_comb \Selector0~36 (
// Equation(s):
// \Selector0~36_combout  = (Mux292 & (((\ShiftLeft0~8_combout ) # (\ShiftLeft0~9_combout )))) # (!Mux292 & (\ShiftLeft0~13_combout ))

	.dataa(Mux292),
	.datab(\ShiftLeft0~13_combout ),
	.datac(\ShiftLeft0~8_combout ),
	.datad(\ShiftLeft0~9_combout ),
	.cin(gnd),
	.combout(\Selector0~36_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~36 .lut_mask = 16'hEEE4;
defparam \Selector0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N18
cycloneive_lcell_comb \Selector1~9 (
// Equation(s):
// \Selector1~9_combout  = (cuifALUOP_3) # ((!\ShiftRight0~22_combout  & ((Mux28) # (Mux272))))

	.dataa(Mux28),
	.datab(cuifALUOP_3),
	.datac(Mux272),
	.datad(\ShiftRight0~22_combout ),
	.cin(gnd),
	.combout(\Selector1~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~9 .lut_mask = 16'hCCFE;
defparam \Selector1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N16
cycloneive_lcell_comb \Selector16~0 (
// Equation(s):
// \Selector16~0_combout  = (!cuifALUOP_1 & (!\ShiftRight0~22_combout  & (!cuifALUOP_2 & !\Selector1~9_combout )))

	.dataa(cuifALUOP_1),
	.datab(\ShiftRight0~22_combout ),
	.datac(cuifALUOP_2),
	.datad(\Selector1~9_combout ),
	.cin(gnd),
	.combout(\Selector16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~0 .lut_mask = 16'h0001;
defparam \Selector16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N2
cycloneive_lcell_comb \Selector0~23 (
// Equation(s):
// \Selector0~23_combout  = (!cuifALUOP_0 & \Selector16~0_combout )

	.dataa(cuifALUOP_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\Selector16~0_combout ),
	.cin(gnd),
	.combout(\Selector0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~23 .lut_mask = 16'h5500;
defparam \Selector0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N16
cycloneive_lcell_comb \Selector1~10 (
// Equation(s):
// \Selector1~10_combout  = (Mux292) # ((!Mux302 & Mux312))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(gnd),
	.datad(Mux292),
	.cin(gnd),
	.combout(\Selector1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~10 .lut_mask = 16'hFF44;
defparam \Selector1~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N14
cycloneive_lcell_comb \ShiftLeft0~15 (
// Equation(s):
// \ShiftLeft0~15_combout  = (Mux302 & ((Mux312 & (\portB~17_combout )) # (!Mux312 & ((\portB~15_combout )))))

	.dataa(Mux302),
	.datab(portB7),
	.datac(Mux312),
	.datad(portB6),
	.cin(gnd),
	.combout(\ShiftLeft0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~15 .lut_mask = 16'h8A80;
defparam \ShiftLeft0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N16
cycloneive_lcell_comb \ShiftLeft0~16 (
// Equation(s):
// \ShiftLeft0~16_combout  = (Mux312 & (\portB~13_combout )) # (!Mux312 & ((\portB~11_combout )))

	.dataa(gnd),
	.datab(Mux312),
	.datac(portB5),
	.datad(portB4),
	.cin(gnd),
	.combout(\ShiftLeft0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~16 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N18
cycloneive_lcell_comb \ShiftLeft0~17 (
// Equation(s):
// \ShiftLeft0~17_combout  = (\ShiftLeft0~15_combout ) # ((!Mux302 & \ShiftLeft0~16_combout ))

	.dataa(Mux302),
	.datab(gnd),
	.datac(\ShiftLeft0~15_combout ),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~17 .lut_mask = 16'hF5F0;
defparam \ShiftLeft0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N20
cycloneive_lcell_comb \Selector0~25 (
// Equation(s):
// \Selector0~25_combout  = (\Selector0~24_combout  & (((\ShiftLeft0~17_combout ) # (!\Selector1~10_combout )))) # (!\Selector0~24_combout  & (\portB~5_combout  & (\Selector1~10_combout )))

	.dataa(\Selector0~24_combout ),
	.datab(portB1),
	.datac(\Selector1~10_combout ),
	.datad(\ShiftLeft0~17_combout ),
	.cin(gnd),
	.combout(\Selector0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~25 .lut_mask = 16'hEA4A;
defparam \Selector0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N8
cycloneive_lcell_comb \Selector0~26 (
// Equation(s):
// \Selector0~26_combout  = (\Selector0~22_combout  & ((\Selector0~36_combout ) # ((\Selector0~23_combout  & \Selector0~25_combout )))) # (!\Selector0~22_combout  & (((\Selector0~23_combout  & \Selector0~25_combout ))))

	.dataa(\Selector0~22_combout ),
	.datab(\Selector0~36_combout ),
	.datac(\Selector0~23_combout ),
	.datad(\Selector0~25_combout ),
	.cin(gnd),
	.combout(\Selector0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~26 .lut_mask = 16'hF888;
defparam \Selector0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N4
cycloneive_lcell_comb \Selector0~21 (
// Equation(s):
// \Selector0~21_combout  = (\portB~3_combout  & ((\Selector0~19_combout ) # ((!\ShiftRight0~23_combout  & Selector8))))

	.dataa(\Selector0~19_combout ),
	.datab(\ShiftRight0~23_combout ),
	.datac(portB),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Selector0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~21 .lut_mask = 16'hB0A0;
defparam \Selector0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N26
cycloneive_lcell_comb \Selector0~29 (
// Equation(s):
// \Selector0~29_combout  = (\Selector0~28_combout ) # ((\Selector0~16_combout ) # ((\Selector0~26_combout ) # (\Selector0~21_combout )))

	.dataa(\Selector0~28_combout ),
	.datab(\Selector0~16_combout ),
	.datac(\Selector0~26_combout ),
	.datad(\Selector0~21_combout ),
	.cin(gnd),
	.combout(\Selector0~29_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~29 .lut_mask = 16'hFFFE;
defparam \Selector0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N12
cycloneive_lcell_comb \Selector0~31 (
// Equation(s):
// \Selector0~31_combout  = (!cuifALUOP_2 & (cuifALUOP_1 & (!cuifALUOP_0 & !cuifALUOP_3)))

	.dataa(cuifALUOP_2),
	.datab(cuifALUOP_1),
	.datac(cuifALUOP_0),
	.datad(cuifALUOP_3),
	.cin(gnd),
	.combout(\Selector0~31_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~31 .lut_mask = 16'h0004;
defparam \Selector0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N4
cycloneive_lcell_comb \Add0~4 (
// Equation(s):
// \Add0~4_combout  = ((\portB~61_combout  $ (Mux292 $ (!\Add0~3 )))) # (GND)
// \Add0~5  = CARRY((\portB~61_combout  & ((Mux292) # (!\Add0~3 ))) # (!\portB~61_combout  & (Mux292 & !\Add0~3 )))

	.dataa(portB29),
	.datab(Mux292),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
// synopsys translate_off
defparam \Add0~4 .lut_mask = 16'h698E;
defparam \Add0~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N6
cycloneive_lcell_comb \Add0~6 (
// Equation(s):
// \Add0~6_combout  = (Mux28 & ((\portB~59_combout  & (\Add0~5  & VCC)) # (!\portB~59_combout  & (!\Add0~5 )))) # (!Mux28 & ((\portB~59_combout  & (!\Add0~5 )) # (!\portB~59_combout  & ((\Add0~5 ) # (GND)))))
// \Add0~7  = CARRY((Mux28 & (!\portB~59_combout  & !\Add0~5 )) # (!Mux28 & ((!\Add0~5 ) # (!\portB~59_combout ))))

	.dataa(Mux28),
	.datab(portB28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
// synopsys translate_off
defparam \Add0~6 .lut_mask = 16'h9617;
defparam \Add0~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N8
cycloneive_lcell_comb \Add0~8 (
// Equation(s):
// \Add0~8_combout  = ((\portB~57_combout  $ (Mux272 $ (!\Add0~7 )))) # (GND)
// \Add0~9  = CARRY((\portB~57_combout  & ((Mux272) # (!\Add0~7 ))) # (!\portB~57_combout  & (Mux272 & !\Add0~7 )))

	.dataa(portB27),
	.datab(Mux272),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
// synopsys translate_off
defparam \Add0~8 .lut_mask = 16'h698E;
defparam \Add0~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N10
cycloneive_lcell_comb \Add0~10 (
// Equation(s):
// \Add0~10_combout  = (Mux26 & ((\portB~55_combout  & (\Add0~9  & VCC)) # (!\portB~55_combout  & (!\Add0~9 )))) # (!Mux26 & ((\portB~55_combout  & (!\Add0~9 )) # (!\portB~55_combout  & ((\Add0~9 ) # (GND)))))
// \Add0~11  = CARRY((Mux26 & (!\portB~55_combout  & !\Add0~9 )) # (!Mux26 & ((!\Add0~9 ) # (!\portB~55_combout ))))

	.dataa(Mux26),
	.datab(portB26),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
// synopsys translate_off
defparam \Add0~10 .lut_mask = 16'h9617;
defparam \Add0~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N12
cycloneive_lcell_comb \Add0~12 (
// Equation(s):
// \Add0~12_combout  = ((Mux252 $ (\portB~53_combout  $ (!\Add0~11 )))) # (GND)
// \Add0~13  = CARRY((Mux252 & ((\portB~53_combout ) # (!\Add0~11 ))) # (!Mux252 & (\portB~53_combout  & !\Add0~11 )))

	.dataa(Mux252),
	.datab(portB25),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
// synopsys translate_off
defparam \Add0~12 .lut_mask = 16'h698E;
defparam \Add0~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N14
cycloneive_lcell_comb \Add0~14 (
// Equation(s):
// \Add0~14_combout  = (Mux242 & ((\portB~51_combout  & (\Add0~13  & VCC)) # (!\portB~51_combout  & (!\Add0~13 )))) # (!Mux242 & ((\portB~51_combout  & (!\Add0~13 )) # (!\portB~51_combout  & ((\Add0~13 ) # (GND)))))
// \Add0~15  = CARRY((Mux242 & (!\portB~51_combout  & !\Add0~13 )) # (!Mux242 & ((!\Add0~13 ) # (!\portB~51_combout ))))

	.dataa(Mux242),
	.datab(portB24),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
// synopsys translate_off
defparam \Add0~14 .lut_mask = 16'h9617;
defparam \Add0~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N16
cycloneive_lcell_comb \Add0~16 (
// Equation(s):
// \Add0~16_combout  = ((\portB~49_combout  $ (Mux23 $ (!\Add0~15 )))) # (GND)
// \Add0~17  = CARRY((\portB~49_combout  & ((Mux23) # (!\Add0~15 ))) # (!\portB~49_combout  & (Mux23 & !\Add0~15 )))

	.dataa(portB23),
	.datab(Mux23),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
// synopsys translate_off
defparam \Add0~16 .lut_mask = 16'h698E;
defparam \Add0~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N18
cycloneive_lcell_comb \Add0~18 (
// Equation(s):
// \Add0~18_combout  = (Mux22 & ((\portB~47_combout  & (\Add0~17  & VCC)) # (!\portB~47_combout  & (!\Add0~17 )))) # (!Mux22 & ((\portB~47_combout  & (!\Add0~17 )) # (!\portB~47_combout  & ((\Add0~17 ) # (GND)))))
// \Add0~19  = CARRY((Mux22 & (!\portB~47_combout  & !\Add0~17 )) # (!Mux22 & ((!\Add0~17 ) # (!\portB~47_combout ))))

	.dataa(Mux22),
	.datab(portB22),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
// synopsys translate_off
defparam \Add0~18 .lut_mask = 16'h9617;
defparam \Add0~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N20
cycloneive_lcell_comb \Add0~20 (
// Equation(s):
// \Add0~20_combout  = ((Mux21 $ (\portB~45_combout  $ (!\Add0~19 )))) # (GND)
// \Add0~21  = CARRY((Mux21 & ((\portB~45_combout ) # (!\Add0~19 ))) # (!Mux21 & (\portB~45_combout  & !\Add0~19 )))

	.dataa(Mux21),
	.datab(portB21),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
// synopsys translate_off
defparam \Add0~20 .lut_mask = 16'h698E;
defparam \Add0~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N22
cycloneive_lcell_comb \Add0~22 (
// Equation(s):
// \Add0~22_combout  = (\portB~43_combout  & ((Mux20 & (\Add0~21  & VCC)) # (!Mux20 & (!\Add0~21 )))) # (!\portB~43_combout  & ((Mux20 & (!\Add0~21 )) # (!Mux20 & ((\Add0~21 ) # (GND)))))
// \Add0~23  = CARRY((\portB~43_combout  & (!Mux20 & !\Add0~21 )) # (!\portB~43_combout  & ((!\Add0~21 ) # (!Mux20))))

	.dataa(portB20),
	.datab(Mux20),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
// synopsys translate_off
defparam \Add0~22 .lut_mask = 16'h9617;
defparam \Add0~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N24
cycloneive_lcell_comb \Add0~24 (
// Equation(s):
// \Add0~24_combout  = ((Mux19 $ (\portB~41_combout  $ (!\Add0~23 )))) # (GND)
// \Add0~25  = CARRY((Mux19 & ((\portB~41_combout ) # (!\Add0~23 ))) # (!Mux19 & (\portB~41_combout  & !\Add0~23 )))

	.dataa(Mux19),
	.datab(portB19),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
// synopsys translate_off
defparam \Add0~24 .lut_mask = 16'h698E;
defparam \Add0~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N26
cycloneive_lcell_comb \Add0~26 (
// Equation(s):
// \Add0~26_combout  = (\portB~39_combout  & ((Mux18 & (\Add0~25  & VCC)) # (!Mux18 & (!\Add0~25 )))) # (!\portB~39_combout  & ((Mux18 & (!\Add0~25 )) # (!Mux18 & ((\Add0~25 ) # (GND)))))
// \Add0~27  = CARRY((\portB~39_combout  & (!Mux18 & !\Add0~25 )) # (!\portB~39_combout  & ((!\Add0~25 ) # (!Mux18))))

	.dataa(portB18),
	.datab(Mux18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout(\Add0~27 ));
// synopsys translate_off
defparam \Add0~26 .lut_mask = 16'h9617;
defparam \Add0~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N28
cycloneive_lcell_comb \Add0~28 (
// Equation(s):
// \Add0~28_combout  = ((\portB~37_combout  $ (Mux17 $ (!\Add0~27 )))) # (GND)
// \Add0~29  = CARRY((\portB~37_combout  & ((Mux17) # (!\Add0~27 ))) # (!\portB~37_combout  & (Mux17 & !\Add0~27 )))

	.dataa(portB17),
	.datab(Mux17),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~27 ),
	.combout(\Add0~28_combout ),
	.cout(\Add0~29 ));
// synopsys translate_off
defparam \Add0~28 .lut_mask = 16'h698E;
defparam \Add0~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N30
cycloneive_lcell_comb \Add0~30 (
// Equation(s):
// \Add0~30_combout  = (\portB~35_combout  & ((Mux16 & (\Add0~29  & VCC)) # (!Mux16 & (!\Add0~29 )))) # (!\portB~35_combout  & ((Mux16 & (!\Add0~29 )) # (!Mux16 & ((\Add0~29 ) # (GND)))))
// \Add0~31  = CARRY((\portB~35_combout  & (!Mux16 & !\Add0~29 )) # (!\portB~35_combout  & ((!\Add0~29 ) # (!Mux16))))

	.dataa(portB16),
	.datab(Mux16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~29 ),
	.combout(\Add0~30_combout ),
	.cout(\Add0~31 ));
// synopsys translate_off
defparam \Add0~30 .lut_mask = 16'h9617;
defparam \Add0~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N0
cycloneive_lcell_comb \Add0~32 (
// Equation(s):
// \Add0~32_combout  = ((\portB~33_combout  $ (Mux15 $ (!\Add0~31 )))) # (GND)
// \Add0~33  = CARRY((\portB~33_combout  & ((Mux15) # (!\Add0~31 ))) # (!\portB~33_combout  & (Mux15 & !\Add0~31 )))

	.dataa(portB15),
	.datab(Mux15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~31 ),
	.combout(\Add0~32_combout ),
	.cout(\Add0~33 ));
// synopsys translate_off
defparam \Add0~32 .lut_mask = 16'h698E;
defparam \Add0~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N2
cycloneive_lcell_comb \Add0~34 (
// Equation(s):
// \Add0~34_combout  = (\portB~31_combout  & ((Mux14 & (\Add0~33  & VCC)) # (!Mux14 & (!\Add0~33 )))) # (!\portB~31_combout  & ((Mux14 & (!\Add0~33 )) # (!Mux14 & ((\Add0~33 ) # (GND)))))
// \Add0~35  = CARRY((\portB~31_combout  & (!Mux14 & !\Add0~33 )) # (!\portB~31_combout  & ((!\Add0~33 ) # (!Mux14))))

	.dataa(portB14),
	.datab(Mux14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~33 ),
	.combout(\Add0~34_combout ),
	.cout(\Add0~35 ));
// synopsys translate_off
defparam \Add0~34 .lut_mask = 16'h9617;
defparam \Add0~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N4
cycloneive_lcell_comb \Add0~36 (
// Equation(s):
// \Add0~36_combout  = ((\portB~29_combout  $ (Mux13 $ (!\Add0~35 )))) # (GND)
// \Add0~37  = CARRY((\portB~29_combout  & ((Mux13) # (!\Add0~35 ))) # (!\portB~29_combout  & (Mux13 & !\Add0~35 )))

	.dataa(portB13),
	.datab(Mux13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~35 ),
	.combout(\Add0~36_combout ),
	.cout(\Add0~37 ));
// synopsys translate_off
defparam \Add0~36 .lut_mask = 16'h698E;
defparam \Add0~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N6
cycloneive_lcell_comb \Add0~38 (
// Equation(s):
// \Add0~38_combout  = (\portB~27_combout  & ((Mux12 & (\Add0~37  & VCC)) # (!Mux12 & (!\Add0~37 )))) # (!\portB~27_combout  & ((Mux12 & (!\Add0~37 )) # (!Mux12 & ((\Add0~37 ) # (GND)))))
// \Add0~39  = CARRY((\portB~27_combout  & (!Mux12 & !\Add0~37 )) # (!\portB~27_combout  & ((!\Add0~37 ) # (!Mux12))))

	.dataa(portB12),
	.datab(Mux12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~37 ),
	.combout(\Add0~38_combout ),
	.cout(\Add0~39 ));
// synopsys translate_off
defparam \Add0~38 .lut_mask = 16'h9617;
defparam \Add0~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N8
cycloneive_lcell_comb \Add0~40 (
// Equation(s):
// \Add0~40_combout  = ((Mux11 $ (\portB~25_combout  $ (!\Add0~39 )))) # (GND)
// \Add0~41  = CARRY((Mux11 & ((\portB~25_combout ) # (!\Add0~39 ))) # (!Mux11 & (\portB~25_combout  & !\Add0~39 )))

	.dataa(Mux11),
	.datab(portB11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~39 ),
	.combout(\Add0~40_combout ),
	.cout(\Add0~41 ));
// synopsys translate_off
defparam \Add0~40 .lut_mask = 16'h698E;
defparam \Add0~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N10
cycloneive_lcell_comb \Add0~42 (
// Equation(s):
// \Add0~42_combout  = (Mux10 & ((\portB~23_combout  & (\Add0~41  & VCC)) # (!\portB~23_combout  & (!\Add0~41 )))) # (!Mux10 & ((\portB~23_combout  & (!\Add0~41 )) # (!\portB~23_combout  & ((\Add0~41 ) # (GND)))))
// \Add0~43  = CARRY((Mux10 & (!\portB~23_combout  & !\Add0~41 )) # (!Mux10 & ((!\Add0~41 ) # (!\portB~23_combout ))))

	.dataa(Mux10),
	.datab(portB10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~41 ),
	.combout(\Add0~42_combout ),
	.cout(\Add0~43 ));
// synopsys translate_off
defparam \Add0~42 .lut_mask = 16'h9617;
defparam \Add0~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N12
cycloneive_lcell_comb \Add0~44 (
// Equation(s):
// \Add0~44_combout  = ((Mux9 $ (\portB~21_combout  $ (!\Add0~43 )))) # (GND)
// \Add0~45  = CARRY((Mux9 & ((\portB~21_combout ) # (!\Add0~43 ))) # (!Mux9 & (\portB~21_combout  & !\Add0~43 )))

	.dataa(Mux9),
	.datab(portB9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~43 ),
	.combout(\Add0~44_combout ),
	.cout(\Add0~45 ));
// synopsys translate_off
defparam \Add0~44 .lut_mask = 16'h698E;
defparam \Add0~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N14
cycloneive_lcell_comb \Add0~46 (
// Equation(s):
// \Add0~46_combout  = (\portB~19_combout  & ((Mux8 & (\Add0~45  & VCC)) # (!Mux8 & (!\Add0~45 )))) # (!\portB~19_combout  & ((Mux8 & (!\Add0~45 )) # (!Mux8 & ((\Add0~45 ) # (GND)))))
// \Add0~47  = CARRY((\portB~19_combout  & (!Mux8 & !\Add0~45 )) # (!\portB~19_combout  & ((!\Add0~45 ) # (!Mux8))))

	.dataa(portB8),
	.datab(Mux8),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~45 ),
	.combout(\Add0~46_combout ),
	.cout(\Add0~47 ));
// synopsys translate_off
defparam \Add0~46 .lut_mask = 16'h9617;
defparam \Add0~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N16
cycloneive_lcell_comb \Add0~48 (
// Equation(s):
// \Add0~48_combout  = ((Mux72 $ (\portB~17_combout  $ (!\Add0~47 )))) # (GND)
// \Add0~49  = CARRY((Mux72 & ((\portB~17_combout ) # (!\Add0~47 ))) # (!Mux72 & (\portB~17_combout  & !\Add0~47 )))

	.dataa(Mux72),
	.datab(portB7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~47 ),
	.combout(\Add0~48_combout ),
	.cout(\Add0~49 ));
// synopsys translate_off
defparam \Add0~48 .lut_mask = 16'h698E;
defparam \Add0~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N18
cycloneive_lcell_comb \Add0~50 (
// Equation(s):
// \Add0~50_combout  = (\portB~15_combout  & ((Mux6 & (\Add0~49  & VCC)) # (!Mux6 & (!\Add0~49 )))) # (!\portB~15_combout  & ((Mux6 & (!\Add0~49 )) # (!Mux6 & ((\Add0~49 ) # (GND)))))
// \Add0~51  = CARRY((\portB~15_combout  & (!Mux6 & !\Add0~49 )) # (!\portB~15_combout  & ((!\Add0~49 ) # (!Mux6))))

	.dataa(portB6),
	.datab(Mux6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~49 ),
	.combout(\Add0~50_combout ),
	.cout(\Add0~51 ));
// synopsys translate_off
defparam \Add0~50 .lut_mask = 16'h9617;
defparam \Add0~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N20
cycloneive_lcell_comb \Add0~52 (
// Equation(s):
// \Add0~52_combout  = ((\portB~13_combout  $ (Mux5 $ (!\Add0~51 )))) # (GND)
// \Add0~53  = CARRY((\portB~13_combout  & ((Mux5) # (!\Add0~51 ))) # (!\portB~13_combout  & (Mux5 & !\Add0~51 )))

	.dataa(portB5),
	.datab(Mux5),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~51 ),
	.combout(\Add0~52_combout ),
	.cout(\Add0~53 ));
// synopsys translate_off
defparam \Add0~52 .lut_mask = 16'h698E;
defparam \Add0~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N22
cycloneive_lcell_comb \Add0~54 (
// Equation(s):
// \Add0~54_combout  = (\portB~11_combout  & ((Mux4 & (\Add0~53  & VCC)) # (!Mux4 & (!\Add0~53 )))) # (!\portB~11_combout  & ((Mux4 & (!\Add0~53 )) # (!Mux4 & ((\Add0~53 ) # (GND)))))
// \Add0~55  = CARRY((\portB~11_combout  & (!Mux4 & !\Add0~53 )) # (!\portB~11_combout  & ((!\Add0~53 ) # (!Mux4))))

	.dataa(portB4),
	.datab(Mux4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~53 ),
	.combout(\Add0~54_combout ),
	.cout(\Add0~55 ));
// synopsys translate_off
defparam \Add0~54 .lut_mask = 16'h9617;
defparam \Add0~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N24
cycloneive_lcell_comb \Add0~56 (
// Equation(s):
// \Add0~56_combout  = ((Mux3 $ (\portB~9_combout  $ (!\Add0~55 )))) # (GND)
// \Add0~57  = CARRY((Mux3 & ((\portB~9_combout ) # (!\Add0~55 ))) # (!Mux3 & (\portB~9_combout  & !\Add0~55 )))

	.dataa(Mux3),
	.datab(portB3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~55 ),
	.combout(\Add0~56_combout ),
	.cout(\Add0~57 ));
// synopsys translate_off
defparam \Add0~56 .lut_mask = 16'h698E;
defparam \Add0~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N26
cycloneive_lcell_comb \Add0~58 (
// Equation(s):
// \Add0~58_combout  = (Mux2 & ((\portB~7_combout  & (\Add0~57  & VCC)) # (!\portB~7_combout  & (!\Add0~57 )))) # (!Mux2 & ((\portB~7_combout  & (!\Add0~57 )) # (!\portB~7_combout  & ((\Add0~57 ) # (GND)))))
// \Add0~59  = CARRY((Mux2 & (!\portB~7_combout  & !\Add0~57 )) # (!Mux2 & ((!\Add0~57 ) # (!\portB~7_combout ))))

	.dataa(Mux2),
	.datab(portB2),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~57 ),
	.combout(\Add0~58_combout ),
	.cout(\Add0~59 ));
// synopsys translate_off
defparam \Add0~58 .lut_mask = 16'h9617;
defparam \Add0~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N28
cycloneive_lcell_comb \Add0~60 (
// Equation(s):
// \Add0~60_combout  = ((Mux1 $ (\portB~5_combout  $ (!\Add0~59 )))) # (GND)
// \Add0~61  = CARRY((Mux1 & ((\portB~5_combout ) # (!\Add0~59 ))) # (!Mux1 & (\portB~5_combout  & !\Add0~59 )))

	.dataa(Mux1),
	.datab(portB1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~59 ),
	.combout(\Add0~60_combout ),
	.cout(\Add0~61 ));
// synopsys translate_off
defparam \Add0~60 .lut_mask = 16'h698E;
defparam \Add0~60 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N30
cycloneive_lcell_comb \Add0~62 (
// Equation(s):
// \Add0~62_combout  = Mux0 $ (\Add0~61  $ (\portB~3_combout ))

	.dataa(gnd),
	.datab(Mux0),
	.datac(gnd),
	.datad(portB),
	.cin(\Add0~61 ),
	.combout(\Add0~62_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~62 .lut_mask = 16'hC33C;
defparam \Add0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N16
cycloneive_lcell_comb \ShiftLeft0~22 (
// Equation(s):
// \ShiftLeft0~22_combout  = (\portB~55_combout  & ((\ShiftRight0~122_combout ) # ((\portB~51_combout  & \ShiftRight0~123_combout )))) # (!\portB~55_combout  & (\portB~51_combout  & (\ShiftRight0~123_combout )))

	.dataa(portB26),
	.datab(portB24),
	.datac(\ShiftRight0~123_combout ),
	.datad(\ShiftRight0~122_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~22 .lut_mask = 16'hEAC0;
defparam \ShiftLeft0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N22
cycloneive_lcell_comb \ShiftLeft0~21 (
// Equation(s):
// \ShiftLeft0~21_combout  = (Mux312 & ((Mux302 & ((\portB~57_combout ))) # (!Mux302 & (\portB~53_combout ))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB25),
	.datad(portB27),
	.cin(gnd),
	.combout(\ShiftLeft0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~21 .lut_mask = 16'hA820;
defparam \ShiftLeft0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N8
cycloneive_lcell_comb \ShiftLeft0~18 (
// Equation(s):
// \ShiftLeft0~18_combout  = (!Mux302 & ((Mux312 & ((\portB~61_combout ))) # (!Mux312 & (\portB~59_combout ))))

	.dataa(Mux312),
	.datab(portB28),
	.datac(portB29),
	.datad(Mux302),
	.cin(gnd),
	.combout(\ShiftLeft0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~18 .lut_mask = 16'h00E4;
defparam \ShiftLeft0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N28
cycloneive_lcell_comb \ShiftLeft0~19 (
// Equation(s):
// \ShiftLeft0~19_combout  = (Mux312 & (\portB~65_combout )) # (!Mux312 & ((\portB~63_combout )))

	.dataa(gnd),
	.datab(portB31),
	.datac(Mux312),
	.datad(portB30),
	.cin(gnd),
	.combout(\ShiftLeft0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~19 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N2
cycloneive_lcell_comb \ShiftLeft0~20 (
// Equation(s):
// \ShiftLeft0~20_combout  = (\ShiftLeft0~18_combout ) # ((\ShiftLeft0~19_combout  & Mux302))

	.dataa(gnd),
	.datab(\ShiftLeft0~18_combout ),
	.datac(\ShiftLeft0~19_combout ),
	.datad(Mux302),
	.cin(gnd),
	.combout(\ShiftLeft0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~20 .lut_mask = 16'hFCCC;
defparam \ShiftLeft0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N14
cycloneive_lcell_comb \ShiftLeft0~101 (
// Equation(s):
// \ShiftLeft0~101_combout  = (Mux292 & (((\ShiftLeft0~20_combout )))) # (!Mux292 & ((\ShiftLeft0~22_combout ) # ((\ShiftLeft0~21_combout ))))

	.dataa(Mux292),
	.datab(\ShiftLeft0~22_combout ),
	.datac(\ShiftLeft0~21_combout ),
	.datad(\ShiftLeft0~20_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~101_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~101 .lut_mask = 16'hFE54;
defparam \ShiftLeft0~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N8
cycloneive_lcell_comb \Selector1~8 (
// Equation(s):
// \Selector1~8_combout  = (!cuifALUOP_1 & (!cuifALUOP_3 & (!cuifALUOP_2 & !\ShiftRight0~22_combout )))

	.dataa(cuifALUOP_1),
	.datab(cuifALUOP_3),
	.datac(cuifALUOP_2),
	.datad(\ShiftRight0~22_combout ),
	.cin(gnd),
	.combout(\Selector1~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~8 .lut_mask = 16'h0001;
defparam \Selector1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N12
cycloneive_lcell_comb \Selector1~11 (
// Equation(s):
// \Selector1~11_combout  = (!cuifALUOP_0 & (Mux272 & \Selector1~8_combout ))

	.dataa(cuifALUOP_0),
	.datab(gnd),
	.datac(Mux272),
	.datad(\Selector1~8_combout ),
	.cin(gnd),
	.combout(\Selector1~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~11 .lut_mask = 16'h5000;
defparam \Selector1~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N16
cycloneive_lcell_comb \Selector0~30 (
// Equation(s):
// \Selector0~30_combout  = (\Selector1~11_combout  & ((Mux28 & ((\ShiftLeft0~101_combout ))) # (!Mux28 & (\Selector8~1_combout ))))

	.dataa(\Selector8~1_combout ),
	.datab(\ShiftLeft0~101_combout ),
	.datac(Mux28),
	.datad(\Selector1~11_combout ),
	.cin(gnd),
	.combout(\Selector0~30_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~30 .lut_mask = 16'hCA00;
defparam \Selector0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N16
cycloneive_lcell_comb \Selector0~32 (
// Equation(s):
// \Selector0~32_combout  = (\Selector0~30_combout ) # ((\Selector0~31_combout  & \Add0~62_combout ))

	.dataa(\Selector0~31_combout ),
	.datab(gnd),
	.datac(\Add0~62_combout ),
	.datad(\Selector0~30_combout ),
	.cin(gnd),
	.combout(\Selector0~32_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~32 .lut_mask = 16'hFFA0;
defparam \Selector0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N30
cycloneive_lcell_comb \ShiftRight0~52 (
// Equation(s):
// \ShiftRight0~52_combout  = (Mux312 & (!Mux302 & \portB~51_combout ))

	.dataa(gnd),
	.datab(Mux312),
	.datac(Mux302),
	.datad(portB24),
	.cin(gnd),
	.combout(\ShiftRight0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~52 .lut_mask = 16'h0C00;
defparam \ShiftRight0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N18
cycloneive_lcell_comb \ShiftLeft0~43 (
// Equation(s):
// \ShiftLeft0~43_combout  = (Mux302 & ((Mux312 & ((\portB~55_combout ))) # (!Mux312 & (\portB~53_combout ))))

	.dataa(portB25),
	.datab(Mux312),
	.datac(Mux302),
	.datad(portB26),
	.cin(gnd),
	.combout(\ShiftLeft0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~43 .lut_mask = 16'hE020;
defparam \ShiftLeft0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N8
cycloneive_lcell_comb \ShiftLeft0~44 (
// Equation(s):
// \ShiftLeft0~44_combout  = (\ShiftRight0~52_combout ) # ((\ShiftLeft0~43_combout ) # ((\ShiftRight0~123_combout  & \portB~49_combout )))

	.dataa(\ShiftRight0~123_combout ),
	.datab(portB23),
	.datac(\ShiftRight0~52_combout ),
	.datad(\ShiftLeft0~43_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~44 .lut_mask = 16'hFFF8;
defparam \ShiftLeft0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N20
cycloneive_lcell_comb \ShiftLeft0~45 (
// Equation(s):
// \ShiftLeft0~45_combout  = (Mux312 & ((Mux302 & ((\portB~47_combout ))) # (!Mux302 & (\portB~43_combout ))))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB20),
	.datad(portB22),
	.cin(gnd),
	.combout(\ShiftLeft0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~45 .lut_mask = 16'hC840;
defparam \ShiftLeft0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N30
cycloneive_lcell_comb \Selector11~10 (
// Equation(s):
// \Selector11~10_combout  = (Mux292 & (((\ShiftLeft0~44_combout )))) # (!Mux292 & ((\ShiftLeft0~46_combout ) # ((\ShiftLeft0~45_combout ))))

	.dataa(\ShiftLeft0~46_combout ),
	.datab(Mux292),
	.datac(\ShiftLeft0~44_combout ),
	.datad(\ShiftLeft0~45_combout ),
	.cin(gnd),
	.combout(\Selector11~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~10 .lut_mask = 16'hF3E2;
defparam \Selector11~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N26
cycloneive_lcell_comb \ShiftLeft0~40 (
// Equation(s):
// \ShiftLeft0~40_combout  = (Mux302 & ((Mux312 & (\portB~63_combout )) # (!Mux312 & ((\portB~61_combout )))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB30),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~40 .lut_mask = 16'hC480;
defparam \ShiftLeft0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N16
cycloneive_lcell_comb \ShiftLeft0~41 (
// Equation(s):
// \ShiftLeft0~41_combout  = (\ShiftLeft0~40_combout ) # ((Mux312 & (!Mux302 & \portB~59_combout )))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(\ShiftLeft0~40_combout ),
	.datad(portB28),
	.cin(gnd),
	.combout(\ShiftLeft0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~41 .lut_mask = 16'hF2F0;
defparam \ShiftLeft0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N22
cycloneive_lcell_comb \ShiftLeft0~42 (
// Equation(s):
// \ShiftLeft0~42_combout  = (\ShiftLeft0~41_combout ) # ((\ShiftRight0~123_combout  & \portB~57_combout ))

	.dataa(\ShiftRight0~123_combout ),
	.datab(gnd),
	.datac(portB27),
	.datad(\ShiftLeft0~41_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~42 .lut_mask = 16'hFFA0;
defparam \ShiftLeft0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N12
cycloneive_lcell_comb \ShiftLeft0~102 (
// Equation(s):
// \ShiftLeft0~102_combout  = (Mux292 & (\portB~65_combout  & (\ShiftRight0~123_combout ))) # (!Mux292 & (((\ShiftLeft0~42_combout ))))

	.dataa(portB31),
	.datab(Mux292),
	.datac(\ShiftRight0~123_combout ),
	.datad(\ShiftLeft0~42_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~102_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~102 .lut_mask = 16'hB380;
defparam \ShiftLeft0~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N6
cycloneive_lcell_comb \ShiftLeft0~48 (
// Equation(s):
// \ShiftLeft0~48_combout  = (Mux28 & ((\ShiftLeft0~102_combout ))) # (!Mux28 & (\Selector11~10_combout ))

	.dataa(gnd),
	.datab(Mux28),
	.datac(\Selector11~10_combout ),
	.datad(\ShiftLeft0~102_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~48 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N30
cycloneive_lcell_comb \Selector0~27 (
// Equation(s):
// \Selector0~27_combout  = (cuifALUOP_0 & (cuifALUOP_1 & (!cuifALUOP_3 & cuifALUOP_2)))

	.dataa(cuifALUOP_0),
	.datab(cuifALUOP_1),
	.datac(cuifALUOP_3),
	.datad(cuifALUOP_2),
	.cin(gnd),
	.combout(\Selector0~27_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~27 .lut_mask = 16'h0800;
defparam \Selector0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N30
cycloneive_lcell_comb \Selector3~1 (
// Equation(s):
// \Selector3~1_combout  = (\portB~9_combout  & (\Selector0~15_combout  & ((!Mux3)))) # (!\portB~9_combout  & ((Mux3 & (\Selector0~15_combout )) # (!Mux3 & ((\Selector0~27_combout )))))

	.dataa(\Selector0~15_combout ),
	.datab(portB3),
	.datac(\Selector0~27_combout ),
	.datad(Mux3),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~1 .lut_mask = 16'h22B8;
defparam \Selector3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N2
cycloneive_lcell_comb \Selector3~0 (
// Equation(s):
// \Selector3~0_combout  = (\Selector0~31_combout  & ((\Add0~56_combout ) # ((\Selector0~14_combout  & \Add1~56_combout )))) # (!\Selector0~31_combout  & (\Selector0~14_combout  & ((\Add1~56_combout ))))

	.dataa(\Selector0~31_combout ),
	.datab(\Selector0~14_combout ),
	.datac(\Add0~56_combout ),
	.datad(\Add1~56_combout ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~0 .lut_mask = 16'hECA0;
defparam \Selector3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N4
cycloneive_lcell_comb \Selector3~2 (
// Equation(s):
// \Selector3~2_combout  = (\Selector3~1_combout ) # ((\Selector3~0_combout ) # ((Mux3 & \Selector0~17_combout )))

	.dataa(Mux3),
	.datab(\Selector0~17_combout ),
	.datac(\Selector3~1_combout ),
	.datad(\Selector3~0_combout ),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~2 .lut_mask = 16'hFFF8;
defparam \Selector3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N16
cycloneive_lcell_comb \ShiftRight0~124 (
// Equation(s):
// \ShiftRight0~124_combout  = (!Mux28 & ((dcifimemload_25 & (!Mux29)) # (!dcifimemload_25 & ((!Mux291)))))

	.dataa(Mux29),
	.datab(dcifimemload_25),
	.datac(Mux291),
	.datad(Mux28),
	.cin(gnd),
	.combout(\ShiftRight0~124_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~124 .lut_mask = 16'h0047;
defparam \ShiftRight0~124 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N22
cycloneive_lcell_comb \Selector3~3 (
// Equation(s):
// \Selector3~3_combout  = (\ShiftRight0~124_combout  & (Selector8 & \ShiftRight0~26_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~124_combout ),
	.datac(Selector8),
	.datad(\ShiftRight0~26_combout ),
	.cin(gnd),
	.combout(\Selector3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~3 .lut_mask = 16'hC000;
defparam \Selector3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N22
cycloneive_lcell_comb \Selector0~18 (
// Equation(s):
// \Selector0~18_combout  = (!cuifALUOP_3 & (!cuifALUOP_1 & (cuifALUOP_2 & !cuifALUOP_0)))

	.dataa(cuifALUOP_3),
	.datab(cuifALUOP_1),
	.datac(cuifALUOP_2),
	.datad(cuifALUOP_0),
	.cin(gnd),
	.combout(\Selector0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~18 .lut_mask = 16'h0010;
defparam \Selector0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N24
cycloneive_lcell_comb \Selector3~4 (
// Equation(s):
// \Selector3~4_combout  = (\portB~9_combout  & ((\Selector0~17_combout ) # ((Mux3 & \Selector0~18_combout ))))

	.dataa(Mux3),
	.datab(\Selector0~18_combout ),
	.datac(\Selector0~17_combout ),
	.datad(portB3),
	.cin(gnd),
	.combout(\Selector3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~4 .lut_mask = 16'hF800;
defparam \Selector3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N18
cycloneive_lcell_comb \Selector3~5 (
// Equation(s):
// \Selector3~5_combout  = (cuifALUOP_3) # ((cuifALUOP_2) # ((Mux272 & !\ShiftRight0~22_combout )))

	.dataa(cuifALUOP_3),
	.datab(cuifALUOP_2),
	.datac(Mux272),
	.datad(\ShiftRight0~22_combout ),
	.cin(gnd),
	.combout(\Selector3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~5 .lut_mask = 16'hEEFE;
defparam \Selector3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N26
cycloneive_lcell_comb \Selector2~0 (
// Equation(s):
// \Selector2~0_combout  = (!cuifALUOP_0 & (!\ShiftRight0~22_combout  & (!cuifALUOP_1 & !\Selector3~5_combout )))

	.dataa(cuifALUOP_0),
	.datab(\ShiftRight0~22_combout ),
	.datac(cuifALUOP_1),
	.datad(\Selector3~5_combout ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~0 .lut_mask = 16'h0001;
defparam \Selector2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N16
cycloneive_lcell_comb \ShiftLeft0~29 (
// Equation(s):
// \ShiftLeft0~29_combout  = (Mux312 & (\portB~15_combout )) # (!Mux312 & ((\portB~13_combout )))

	.dataa(Mux312),
	.datab(gnd),
	.datac(portB6),
	.datad(portB5),
	.cin(gnd),
	.combout(\ShiftLeft0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~29 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N24
cycloneive_lcell_comb \ShiftLeft0~37 (
// Equation(s):
// \ShiftLeft0~37_combout  = (\portB~33_combout  & ((\ShiftRight0~123_combout ) # ((\portB~37_combout  & \ShiftRight0~122_combout )))) # (!\portB~33_combout  & (\portB~37_combout  & ((\ShiftRight0~122_combout ))))

	.dataa(portB15),
	.datab(portB17),
	.datac(\ShiftRight0~123_combout ),
	.datad(\ShiftRight0~122_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~37 .lut_mask = 16'hECA0;
defparam \ShiftLeft0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N8
cycloneive_lcell_comb \ShiftLeft0~33 (
// Equation(s):
// \ShiftLeft0~33_combout  = (Mux312 & ((Mux302 & (\portB~31_combout )) # (!Mux302 & ((\portB~27_combout )))))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB14),
	.datad(portB12),
	.cin(gnd),
	.combout(\ShiftLeft0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~33 .lut_mask = 16'hC480;
defparam \ShiftLeft0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N4
cycloneive_lcell_comb \ShiftLeft0~34 (
// Equation(s):
// \ShiftLeft0~34_combout  = (\ShiftRight0~123_combout  & ((\portB~25_combout ) # ((\ShiftRight0~122_combout  & \portB~29_combout )))) # (!\ShiftRight0~123_combout  & (\ShiftRight0~122_combout  & ((\portB~29_combout ))))

	.dataa(\ShiftRight0~123_combout ),
	.datab(\ShiftRight0~122_combout ),
	.datac(portB11),
	.datad(portB13),
	.cin(gnd),
	.combout(\ShiftLeft0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~34 .lut_mask = 16'hECA0;
defparam \ShiftLeft0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N14
cycloneive_lcell_comb \ShiftLeft0~35 (
// Equation(s):
// \ShiftLeft0~35_combout  = (\ShiftLeft0~33_combout ) # (\ShiftLeft0~34_combout )

	.dataa(gnd),
	.datab(\ShiftLeft0~33_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~34_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~35 .lut_mask = 16'hFFCC;
defparam \ShiftLeft0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N24
cycloneive_lcell_comb \ShiftLeft0~38 (
// Equation(s):
// \ShiftLeft0~38_combout  = (Mux292 & ((\ShiftLeft0~36_combout ) # ((\ShiftLeft0~37_combout )))) # (!Mux292 & (((\ShiftLeft0~35_combout ))))

	.dataa(\ShiftLeft0~36_combout ),
	.datab(Mux292),
	.datac(\ShiftLeft0~37_combout ),
	.datad(\ShiftLeft0~35_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~38 .lut_mask = 16'hFBC8;
defparam \ShiftLeft0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N14
cycloneive_lcell_comb \Selector3~6 (
// Equation(s):
// \Selector3~6_combout  = (Mux28) # ((Mux302 & !Mux292))

	.dataa(gnd),
	.datab(Mux302),
	.datac(Mux292),
	.datad(Mux28),
	.cin(gnd),
	.combout(\Selector3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~6 .lut_mask = 16'hFF0C;
defparam \Selector3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N22
cycloneive_lcell_comb \ShiftRight0~51 (
// Equation(s):
// \ShiftRight0~51_combout  = (!Mux302 & (Mux312 & \portB~19_combout ))

	.dataa(Mux302),
	.datab(gnd),
	.datac(Mux312),
	.datad(portB8),
	.cin(gnd),
	.combout(\ShiftRight0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~51 .lut_mask = 16'h5000;
defparam \ShiftRight0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N20
cycloneive_lcell_comb \ShiftLeft0~30 (
// Equation(s):
// \ShiftLeft0~30_combout  = (Mux302 & ((Mux312 & (\portB~23_combout )) # (!Mux312 & ((\portB~21_combout )))))

	.dataa(Mux302),
	.datab(portB10),
	.datac(portB9),
	.datad(Mux312),
	.cin(gnd),
	.combout(\ShiftLeft0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~30 .lut_mask = 16'h88A0;
defparam \ShiftLeft0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N30
cycloneive_lcell_comb \ShiftLeft0~31 (
// Equation(s):
// \ShiftLeft0~31_combout  = (\ShiftRight0~51_combout ) # ((\ShiftLeft0~30_combout ) # ((\portB~17_combout  & \ShiftRight0~123_combout )))

	.dataa(portB7),
	.datab(\ShiftRight0~123_combout ),
	.datac(\ShiftRight0~51_combout ),
	.datad(\ShiftLeft0~30_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~31 .lut_mask = 16'hFFF8;
defparam \ShiftLeft0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N20
cycloneive_lcell_comb \Selector3~7 (
// Equation(s):
// \Selector3~7_combout  = (\ShiftRight0~124_combout  & (\ShiftLeft0~32_combout  & (!\Selector3~6_combout ))) # (!\ShiftRight0~124_combout  & (((\Selector3~6_combout ) # (\ShiftLeft0~31_combout ))))

	.dataa(\ShiftLeft0~32_combout ),
	.datab(\ShiftRight0~124_combout ),
	.datac(\Selector3~6_combout ),
	.datad(\ShiftLeft0~31_combout ),
	.cin(gnd),
	.combout(\Selector3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~7 .lut_mask = 16'h3B38;
defparam \Selector3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N18
cycloneive_lcell_comb \Selector3~8 (
// Equation(s):
// \Selector3~8_combout  = (\Selector3~6_combout  & ((\Selector3~7_combout  & ((\ShiftLeft0~38_combout ))) # (!\Selector3~7_combout  & (\ShiftLeft0~29_combout )))) # (!\Selector3~6_combout  & (((\Selector3~7_combout ))))

	.dataa(\Selector3~6_combout ),
	.datab(\ShiftLeft0~29_combout ),
	.datac(\ShiftLeft0~38_combout ),
	.datad(\Selector3~7_combout ),
	.cin(gnd),
	.combout(\Selector3~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~8 .lut_mask = 16'hF588;
defparam \Selector3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N16
cycloneive_lcell_comb \Selector3~9 (
// Equation(s):
// \Selector3~9_combout  = (\Selector3~3_combout ) # ((\Selector3~4_combout ) # ((\Selector2~0_combout  & \Selector3~8_combout )))

	.dataa(\Selector3~3_combout ),
	.datab(\Selector3~4_combout ),
	.datac(\Selector2~0_combout ),
	.datad(\Selector3~8_combout ),
	.cin(gnd),
	.combout(\Selector3~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~9 .lut_mask = 16'hFEEE;
defparam \Selector3~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N24
cycloneive_lcell_comb \Selector7~14 (
// Equation(s):
// \Selector7~14_combout  = (\portB~17_combout  & ((\Selector0~5_combout ) # ((Mux72 & \Selector0~6_combout ))))

	.dataa(portB7),
	.datab(Mux72),
	.datac(\Selector0~5_combout ),
	.datad(\Selector0~6_combout ),
	.cin(gnd),
	.combout(\Selector7~14_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~14 .lut_mask = 16'hA8A0;
defparam \Selector7~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N22
cycloneive_lcell_comb \Selector7~15 (
// Equation(s):
// \Selector7~15_combout  = (\Selector7~14_combout ) # ((\Selector0~7_combout  & (!\portB~17_combout  & !Mux72)))

	.dataa(\Selector0~7_combout ),
	.datab(\Selector7~14_combout ),
	.datac(portB7),
	.datad(Mux72),
	.cin(gnd),
	.combout(\Selector7~15_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~15 .lut_mask = 16'hCCCE;
defparam \Selector7~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N4
cycloneive_lcell_comb \Selector7~16 (
// Equation(s):
// \Selector7~16_combout  = (\Selector7~15_combout ) # ((\Selector0~11_combout  & (\portB~17_combout  $ (Mux72))))

	.dataa(portB7),
	.datab(\Selector0~11_combout ),
	.datac(\Selector7~15_combout ),
	.datad(Mux72),
	.cin(gnd),
	.combout(\Selector7~16_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~16 .lut_mask = 16'hF4F8;
defparam \Selector7~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N28
cycloneive_lcell_comb \Selector4~0 (
// Equation(s):
// \Selector4~0_combout  = (!\ShiftRight0~22_combout  & \Selector0~9_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftRight0~22_combout ),
	.datad(\Selector0~9_combout ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~0 .lut_mask = 16'h0F00;
defparam \Selector4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N22
cycloneive_lcell_comb \Selector7~8 (
// Equation(s):
// \Selector7~8_combout  = (\Selector0~5_combout  & ((dcifimemload_25 & ((Mux7))) # (!dcifimemload_25 & (Mux71))))

	.dataa(Mux71),
	.datab(dcifimemload_25),
	.datac(\Selector0~5_combout ),
	.datad(Mux7),
	.cin(gnd),
	.combout(\Selector7~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~8 .lut_mask = 16'hE020;
defparam \Selector7~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N20
cycloneive_lcell_comb \Selector7~10 (
// Equation(s):
// \Selector7~10_combout  = (Mux272) # ((!Mux28 & Mux292))

	.dataa(Mux28),
	.datab(gnd),
	.datac(Mux292),
	.datad(Mux272),
	.cin(gnd),
	.combout(\Selector7~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~10 .lut_mask = 16'hFF50;
defparam \Selector7~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N12
cycloneive_lcell_comb \Selector7~18 (
// Equation(s):
// \Selector7~18_combout  = (Mux28) # ((dcifimemload_25 & (Mux27)) # (!dcifimemload_25 & ((Mux271))))

	.dataa(Mux27),
	.datab(Mux271),
	.datac(dcifimemload_25),
	.datad(Mux28),
	.cin(gnd),
	.combout(\Selector7~18_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~18 .lut_mask = 16'hFFAC;
defparam \Selector7~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N20
cycloneive_lcell_comb \ShiftLeft0~46 (
// Equation(s):
// \ShiftLeft0~46_combout  = (\portB~41_combout  & ((\ShiftRight0~123_combout ) # ((\ShiftRight0~122_combout  & \portB~45_combout )))) # (!\portB~41_combout  & (((\ShiftRight0~122_combout  & \portB~45_combout ))))

	.dataa(portB19),
	.datab(\ShiftRight0~123_combout ),
	.datac(\ShiftRight0~122_combout ),
	.datad(portB21),
	.cin(gnd),
	.combout(\ShiftLeft0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~46 .lut_mask = 16'hF888;
defparam \ShiftLeft0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N2
cycloneive_lcell_comb \ShiftLeft0~47 (
// Equation(s):
// \ShiftLeft0~47_combout  = (\ShiftLeft0~45_combout ) # (\ShiftLeft0~46_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftLeft0~45_combout ),
	.datad(\ShiftLeft0~46_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~47 .lut_mask = 16'hFFF0;
defparam \ShiftLeft0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N18
cycloneive_lcell_comb \ShiftLeft0~49 (
// Equation(s):
// \ShiftLeft0~49_combout  = (Mux292 & (((\ShiftLeft0~47_combout )))) # (!Mux292 & ((\ShiftLeft0~36_combout ) # ((\ShiftLeft0~37_combout ))))

	.dataa(\ShiftLeft0~36_combout ),
	.datab(Mux292),
	.datac(\ShiftLeft0~37_combout ),
	.datad(\ShiftLeft0~47_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~49 .lut_mask = 16'hFE32;
defparam \ShiftLeft0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N8
cycloneive_lcell_comb \Selector7~11 (
// Equation(s):
// \Selector7~11_combout  = (\Selector7~10_combout  & (\Selector7~18_combout )) # (!\Selector7~10_combout  & ((\Selector7~18_combout  & ((\ShiftLeft0~49_combout ))) # (!\Selector7~18_combout  & (\ShiftLeft0~31_combout ))))

	.dataa(\Selector7~10_combout ),
	.datab(\Selector7~18_combout ),
	.datac(\ShiftLeft0~31_combout ),
	.datad(\ShiftLeft0~49_combout ),
	.cin(gnd),
	.combout(\Selector7~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~11 .lut_mask = 16'hDC98;
defparam \Selector7~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N30
cycloneive_lcell_comb \ShiftLeft0~39 (
// Equation(s):
// \ShiftLeft0~39_combout  = (\ShiftRight0~123_combout  & \portB~65_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftRight0~123_combout ),
	.datad(portB31),
	.cin(gnd),
	.combout(\ShiftLeft0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~39 .lut_mask = 16'hF000;
defparam \ShiftLeft0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N28
cycloneive_lcell_comb \ShiftLeft0~50 (
// Equation(s):
// \ShiftLeft0~50_combout  = (Mux292 & (!Mux28 & (\ShiftLeft0~42_combout ))) # (!Mux292 & (Mux28 & ((\ShiftLeft0~39_combout ))))

	.dataa(Mux292),
	.datab(Mux28),
	.datac(\ShiftLeft0~42_combout ),
	.datad(\ShiftLeft0~39_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~50_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~50 .lut_mask = 16'h6420;
defparam \ShiftLeft0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N14
cycloneive_lcell_comb \ShiftLeft0~51 (
// Equation(s):
// \ShiftLeft0~51_combout  = (\ShiftLeft0~50_combout ) # ((\ShiftLeft0~44_combout  & \ShiftRight0~124_combout ))

	.dataa(\ShiftLeft0~44_combout ),
	.datab(\ShiftRight0~124_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~50_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~51 .lut_mask = 16'hFF88;
defparam \ShiftLeft0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N22
cycloneive_lcell_comb \Selector7~12 (
// Equation(s):
// \Selector7~12_combout  = (\Selector7~10_combout  & ((\Selector7~11_combout  & ((\ShiftLeft0~51_combout ))) # (!\Selector7~11_combout  & (\ShiftLeft0~35_combout )))) # (!\Selector7~10_combout  & (((\Selector7~11_combout ))))

	.dataa(\ShiftLeft0~35_combout ),
	.datab(\Selector7~10_combout ),
	.datac(\Selector7~11_combout ),
	.datad(\ShiftLeft0~51_combout ),
	.cin(gnd),
	.combout(\Selector7~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~12 .lut_mask = 16'hF838;
defparam \Selector7~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N20
cycloneive_lcell_comb \Selector7~9 (
// Equation(s):
// \Selector7~9_combout  = (\Selector0~10_combout  & ((\Add0~48_combout ) # ((\Selector0~8_combout  & \Add1~48_combout )))) # (!\Selector0~10_combout  & (\Selector0~8_combout  & (\Add1~48_combout )))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~8_combout ),
	.datac(\Add1~48_combout ),
	.datad(\Add0~48_combout ),
	.cin(gnd),
	.combout(\Selector7~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~9 .lut_mask = 16'hEAC0;
defparam \Selector7~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N16
cycloneive_lcell_comb \Selector7~13 (
// Equation(s):
// \Selector7~13_combout  = (\Selector7~8_combout ) # ((\Selector7~9_combout ) # ((\Selector4~0_combout  & \Selector7~12_combout )))

	.dataa(\Selector4~0_combout ),
	.datab(\Selector7~8_combout ),
	.datac(\Selector7~12_combout ),
	.datad(\Selector7~9_combout ),
	.cin(gnd),
	.combout(\Selector7~13_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~13 .lut_mask = 16'hFFEC;
defparam \Selector7~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N20
cycloneive_lcell_comb \Selector0~22 (
// Equation(s):
// \Selector0~22_combout  = (!Mux272 & (Mux28 & (\Selector1~8_combout  & !cuifALUOP_0)))

	.dataa(Mux272),
	.datab(Mux28),
	.datac(\Selector1~8_combout ),
	.datad(cuifALUOP_0),
	.cin(gnd),
	.combout(\Selector0~22_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~22 .lut_mask = 16'h0040;
defparam \Selector0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N28
cycloneive_lcell_comb \Selector8~2 (
// Equation(s):
// \Selector8~2_combout  = (Mux272 & (!Mux28 & (\Selector1~8_combout  & !cuifALUOP_0)))

	.dataa(Mux272),
	.datab(Mux28),
	.datac(\Selector1~8_combout ),
	.datad(cuifALUOP_0),
	.cin(gnd),
	.combout(\Selector8~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~2 .lut_mask = 16'h0020;
defparam \Selector8~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N14
cycloneive_lcell_comb \Selector11~2 (
// Equation(s):
// \Selector11~2_combout  = (\ShiftLeft0~102_combout  & ((\Selector8~2_combout ) # ((\Selector0~22_combout  & \Selector11~10_combout )))) # (!\ShiftLeft0~102_combout  & (\Selector0~22_combout  & (\Selector11~10_combout )))

	.dataa(\ShiftLeft0~102_combout ),
	.datab(\Selector0~22_combout ),
	.datac(\Selector11~10_combout ),
	.datad(\Selector8~2_combout ),
	.cin(gnd),
	.combout(\Selector11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~2 .lut_mask = 16'hEAC0;
defparam \Selector11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N2
cycloneive_lcell_comb \Selector11~4 (
// Equation(s):
// \Selector11~4_combout  = (\portB~25_combout  & ((\Selector0~17_combout ) # ((Mux11 & \Selector0~18_combout ))))

	.dataa(Mux11),
	.datab(\Selector0~17_combout ),
	.datac(portB11),
	.datad(\Selector0~18_combout ),
	.cin(gnd),
	.combout(\Selector11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~4 .lut_mask = 16'hE0C0;
defparam \Selector11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N16
cycloneive_lcell_comb \Selector11~5 (
// Equation(s):
// \Selector11~5_combout  = (\Selector11~4_combout ) # ((!Mux11 & (\Selector0~27_combout  & !\portB~25_combout )))

	.dataa(Mux11),
	.datab(\Selector0~27_combout ),
	.datac(portB11),
	.datad(\Selector11~4_combout ),
	.cin(gnd),
	.combout(\Selector11~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~5 .lut_mask = 16'hFF04;
defparam \Selector11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N22
cycloneive_lcell_comb \Selector11~6 (
// Equation(s):
// \Selector11~6_combout  = (\Selector11~5_combout ) # ((\Selector0~15_combout  & (Mux11 $ (\portB~25_combout ))))

	.dataa(Mux11),
	.datab(\Selector0~15_combout ),
	.datac(portB11),
	.datad(\Selector11~5_combout ),
	.cin(gnd),
	.combout(\Selector11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~6 .lut_mask = 16'hFF48;
defparam \Selector11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N24
cycloneive_lcell_comb \Selector11~3 (
// Equation(s):
// \Selector11~3_combout  = (\Selector0~31_combout  & ((\Add0~40_combout ) # ((\Selector0~14_combout  & \Add1~40_combout )))) # (!\Selector0~31_combout  & (\Selector0~14_combout  & (\Add1~40_combout )))

	.dataa(\Selector0~31_combout ),
	.datab(\Selector0~14_combout ),
	.datac(\Add1~40_combout ),
	.datad(\Add0~40_combout ),
	.cin(gnd),
	.combout(\Selector11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~3 .lut_mask = 16'hEAC0;
defparam \Selector11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N0
cycloneive_lcell_comb \Selector11~7 (
// Equation(s):
// \Selector11~7_combout  = (\Selector11~6_combout ) # ((\Selector11~3_combout ) # ((Mux11 & \Selector0~17_combout )))

	.dataa(Mux11),
	.datab(\Selector0~17_combout ),
	.datac(\Selector11~6_combout ),
	.datad(\Selector11~3_combout ),
	.cin(gnd),
	.combout(\Selector11~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~7 .lut_mask = 16'hFFF8;
defparam \Selector11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N10
cycloneive_lcell_comb \Selector7~19 (
// Equation(s):
// \Selector7~19_combout  = (!Mux28 & ((dcifimemload_25 & (Mux29)) # (!dcifimemload_25 & ((Mux291)))))

	.dataa(Mux29),
	.datab(dcifimemload_25),
	.datac(Mux291),
	.datad(Mux28),
	.cin(gnd),
	.combout(\Selector7~19_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~19 .lut_mask = 16'h00B8;
defparam \Selector7~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N6
cycloneive_lcell_comb \ShiftRight0~53 (
// Equation(s):
// \ShiftRight0~53_combout  = (\ShiftRight0~33_combout  & ((\ShiftRight0~124_combout ) # ((\Selector7~19_combout  & \ShiftRight0~29_combout )))) # (!\ShiftRight0~33_combout  & (((\Selector7~19_combout  & \ShiftRight0~29_combout ))))

	.dataa(\ShiftRight0~33_combout ),
	.datab(\ShiftRight0~124_combout ),
	.datac(\Selector7~19_combout ),
	.datad(\ShiftRight0~29_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~53 .lut_mask = 16'hF888;
defparam \ShiftRight0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N12
cycloneive_lcell_comb \Selector15~0 (
// Equation(s):
// \Selector15~0_combout  = (Mux292 & (\ShiftLeft0~42_combout )) # (!Mux292 & ((\ShiftLeft0~44_combout )))

	.dataa(Mux292),
	.datab(gnd),
	.datac(\ShiftLeft0~42_combout ),
	.datad(\ShiftLeft0~44_combout ),
	.cin(gnd),
	.combout(\Selector15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~0 .lut_mask = 16'hF5A0;
defparam \Selector15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N18
cycloneive_lcell_comb \Selector15~1 (
// Equation(s):
// \Selector15~1_combout  = (\Selector15~0_combout  & ((\Selector0~22_combout ) # ((\ShiftLeft0~49_combout  & \Selector0~23_combout )))) # (!\Selector15~0_combout  & (\ShiftLeft0~49_combout  & ((\Selector0~23_combout ))))

	.dataa(\Selector15~0_combout ),
	.datab(\ShiftLeft0~49_combout ),
	.datac(\Selector0~22_combout ),
	.datad(\Selector0~23_combout ),
	.cin(gnd),
	.combout(\Selector15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~1 .lut_mask = 16'hECA0;
defparam \Selector15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N10
cycloneive_lcell_comb \Selector15~3 (
// Equation(s):
// \Selector15~3_combout  = (\portB~33_combout  & ((\Selector0~17_combout ) # ((Mux15 & \Selector0~18_combout ))))

	.dataa(Mux15),
	.datab(\Selector0~18_combout ),
	.datac(portB15),
	.datad(\Selector0~17_combout ),
	.cin(gnd),
	.combout(\Selector15~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~3 .lut_mask = 16'hF080;
defparam \Selector15~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N28
cycloneive_lcell_comb \Selector15~4 (
// Equation(s):
// \Selector15~4_combout  = (\Selector15~3_combout ) # ((!Mux15 & (\Selector0~27_combout  & !\portB~33_combout )))

	.dataa(Mux15),
	.datab(\Selector0~27_combout ),
	.datac(portB15),
	.datad(\Selector15~3_combout ),
	.cin(gnd),
	.combout(\Selector15~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~4 .lut_mask = 16'hFF04;
defparam \Selector15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N30
cycloneive_lcell_comb \Selector15~5 (
// Equation(s):
// \Selector15~5_combout  = (\Selector15~4_combout ) # ((\Selector0~15_combout  & (Mux15 $ (\portB~33_combout ))))

	.dataa(\Selector0~15_combout ),
	.datab(Mux15),
	.datac(portB15),
	.datad(\Selector15~4_combout ),
	.cin(gnd),
	.combout(\Selector15~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~5 .lut_mask = 16'hFF28;
defparam \Selector15~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N0
cycloneive_lcell_comb \Selector15~2 (
// Equation(s):
// \Selector15~2_combout  = (\Selector0~14_combout  & ((\Add1~32_combout ) # ((\Selector0~31_combout  & \Add0~32_combout )))) # (!\Selector0~14_combout  & (\Selector0~31_combout  & (\Add0~32_combout )))

	.dataa(\Selector0~14_combout ),
	.datab(\Selector0~31_combout ),
	.datac(\Add0~32_combout ),
	.datad(\Add1~32_combout ),
	.cin(gnd),
	.combout(\Selector15~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~2 .lut_mask = 16'hEAC0;
defparam \Selector15~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N20
cycloneive_lcell_comb \Selector15~6 (
// Equation(s):
// \Selector15~6_combout  = (\Selector15~5_combout ) # ((\Selector15~2_combout ) # ((Mux15 & \Selector0~17_combout )))

	.dataa(Mux15),
	.datab(\Selector0~17_combout ),
	.datac(\Selector15~5_combout ),
	.datad(\Selector15~2_combout ),
	.cin(gnd),
	.combout(\Selector15~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~6 .lut_mask = 16'hFFF8;
defparam \Selector15~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N6
cycloneive_lcell_comb \Selector15~7 (
// Equation(s):
// \Selector15~7_combout  = (\Selector15~6_combout ) # ((\portB~65_combout  & (\Selector1~11_combout  & !\ShiftRight0~23_combout )))

	.dataa(portB31),
	.datab(\Selector1~11_combout ),
	.datac(\ShiftRight0~23_combout ),
	.datad(\Selector15~6_combout ),
	.cin(gnd),
	.combout(\Selector15~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~7 .lut_mask = 16'hFF08;
defparam \Selector15~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N14
cycloneive_lcell_comb \Selector28~1 (
// Equation(s):
// \Selector28~1_combout  = (Mux28 & (\Selector0~15_combout  & ((!\portB~59_combout )))) # (!Mux28 & ((\portB~59_combout  & (\Selector0~15_combout )) # (!\portB~59_combout  & ((\Selector0~27_combout )))))

	.dataa(Mux28),
	.datab(\Selector0~15_combout ),
	.datac(\Selector0~27_combout ),
	.datad(portB28),
	.cin(gnd),
	.combout(\Selector28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~1 .lut_mask = 16'h44D8;
defparam \Selector28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N20
cycloneive_lcell_comb \Selector28~0 (
// Equation(s):
// \Selector28~0_combout  = (\Selector0~31_combout  & ((\Add0~6_combout ) # ((\Selector0~14_combout  & \Add1~6_combout )))) # (!\Selector0~31_combout  & (\Selector0~14_combout  & (\Add1~6_combout )))

	.dataa(\Selector0~31_combout ),
	.datab(\Selector0~14_combout ),
	.datac(\Add1~6_combout ),
	.datad(\Add0~6_combout ),
	.cin(gnd),
	.combout(\Selector28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~0 .lut_mask = 16'hEAC0;
defparam \Selector28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N8
cycloneive_lcell_comb \Selector28~2 (
// Equation(s):
// \Selector28~2_combout  = (\Selector28~1_combout ) # ((\Selector28~0_combout ) # ((\Selector0~17_combout  & Mux28)))

	.dataa(\Selector0~17_combout ),
	.datab(Mux28),
	.datac(\Selector28~1_combout ),
	.datad(\Selector28~0_combout ),
	.cin(gnd),
	.combout(\Selector28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~2 .lut_mask = 16'hFFF8;
defparam \Selector28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N14
cycloneive_lcell_comb \Selector16~1 (
// Equation(s):
// \Selector16~1_combout  = (\Selector0~34_combout  & (!Mux272 & !\ShiftRight0~22_combout ))

	.dataa(\Selector0~34_combout ),
	.datab(Mux272),
	.datac(gnd),
	.datad(\ShiftRight0~22_combout ),
	.cin(gnd),
	.combout(\Selector16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~1 .lut_mask = 16'h0022;
defparam \Selector16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N6
cycloneive_lcell_comb \Selector28~3 (
// Equation(s):
// \Selector28~3_combout  = (\ShiftRight0~124_combout  & (\ShiftLeft0~20_combout  & \Selector16~1_combout ))

	.dataa(\ShiftRight0~124_combout ),
	.datab(\ShiftLeft0~20_combout ),
	.datac(gnd),
	.datad(\Selector16~1_combout ),
	.cin(gnd),
	.combout(\Selector28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~3 .lut_mask = 16'h8800;
defparam \Selector28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N24
cycloneive_lcell_comb \Selector28~7 (
// Equation(s):
// \Selector28~7_combout  = (!cuifALUOP_1 & (!\ShiftRight0~22_combout  & (cuifALUOP_0 & !\Selector3~5_combout )))

	.dataa(cuifALUOP_1),
	.datab(\ShiftRight0~22_combout ),
	.datac(cuifALUOP_0),
	.datad(\Selector3~5_combout ),
	.cin(gnd),
	.combout(\Selector28~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~7 .lut_mask = 16'h0010;
defparam \Selector28~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N10
cycloneive_lcell_comb \Selector28~4 (
// Equation(s):
// \Selector28~4_combout  = (\portB~59_combout  & ((\Selector0~17_combout ) # ((Mux28 & \Selector0~18_combout ))))

	.dataa(Mux28),
	.datab(\Selector0~18_combout ),
	.datac(portB28),
	.datad(\Selector0~17_combout ),
	.cin(gnd),
	.combout(\Selector28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~4 .lut_mask = 16'hF080;
defparam \Selector28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N6
cycloneive_lcell_comb \ShiftRight0~55 (
// Equation(s):
// \ShiftRight0~55_combout  = (Mux312 & ((\portB~53_combout ))) # (!Mux312 & (\portB~55_combout ))

	.dataa(portB26),
	.datab(gnd),
	.datac(Mux312),
	.datad(portB25),
	.cin(gnd),
	.combout(\ShiftRight0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~55 .lut_mask = 16'hFA0A;
defparam \ShiftRight0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N14
cycloneive_lcell_comb \ShiftRight0~62 (
// Equation(s):
// \ShiftRight0~62_combout  = (!Mux302 & ((Mux312 & (\portB~41_combout )) # (!Mux312 & ((\portB~43_combout )))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB19),
	.datad(portB20),
	.cin(gnd),
	.combout(\ShiftRight0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~62 .lut_mask = 16'h3120;
defparam \ShiftRight0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N6
cycloneive_lcell_comb \ShiftRight0~60 (
// Equation(s):
// \ShiftRight0~60_combout  = (Mux302 & ((Mux312 & (\portB~29_combout )) # (!Mux312 & ((\portB~31_combout ))))) # (!Mux302 & (((Mux312))))

	.dataa(portB13),
	.datab(Mux302),
	.datac(Mux312),
	.datad(portB14),
	.cin(gnd),
	.combout(\ShiftRight0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~60 .lut_mask = 16'hBCB0;
defparam \ShiftRight0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N8
cycloneive_lcell_comb \ShiftRight0~61 (
// Equation(s):
// \ShiftRight0~61_combout  = (Mux302 & (((\ShiftRight0~60_combout )))) # (!Mux302 & ((\ShiftRight0~60_combout  & (\portB~33_combout )) # (!\ShiftRight0~60_combout  & ((\portB~35_combout )))))

	.dataa(portB15),
	.datab(Mux302),
	.datac(portB16),
	.datad(\ShiftRight0~60_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~61 .lut_mask = 16'hEE30;
defparam \ShiftRight0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N20
cycloneive_lcell_comb \ShiftRight0~63 (
// Equation(s):
// \ShiftRight0~63_combout  = (Mux302 & ((Mux312 & (\portB~37_combout )) # (!Mux312 & ((\portB~39_combout )))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB17),
	.datad(portB18),
	.cin(gnd),
	.combout(\ShiftRight0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~63 .lut_mask = 16'hC480;
defparam \ShiftRight0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N22
cycloneive_lcell_comb \ShiftRight0~64 (
// Equation(s):
// \ShiftRight0~64_combout  = (Mux292 & (((\ShiftRight0~61_combout )))) # (!Mux292 & ((\ShiftRight0~62_combout ) # ((\ShiftRight0~63_combout ))))

	.dataa(Mux292),
	.datab(\ShiftRight0~62_combout ),
	.datac(\ShiftRight0~61_combout ),
	.datad(\ShiftRight0~63_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~64 .lut_mask = 16'hF5E4;
defparam \ShiftRight0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N14
cycloneive_lcell_comb \ShiftRight0~59 (
// Equation(s):
// \ShiftRight0~59_combout  = (Mux312 & ((\portB~57_combout ))) # (!Mux312 & (\portB~59_combout ))

	.dataa(gnd),
	.datab(portB28),
	.datac(portB27),
	.datad(Mux312),
	.cin(gnd),
	.combout(\ShiftRight0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~59 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N10
cycloneive_lcell_comb \ShiftRight0~57 (
// Equation(s):
// \ShiftRight0~57_combout  = (Mux312 & (Mux302 & ((\portB~45_combout )))) # (!Mux312 & (!Mux302 & (\portB~51_combout )))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB24),
	.datad(portB21),
	.cin(gnd),
	.combout(\ShiftRight0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~57 .lut_mask = 16'h9810;
defparam \ShiftRight0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N0
cycloneive_lcell_comb \ShiftRight0~58 (
// Equation(s):
// \ShiftRight0~58_combout  = (\ShiftRight0~56_combout ) # ((\ShiftRight0~57_combout ) # ((\portB~47_combout  & \ShiftRight0~122_combout )))

	.dataa(\ShiftRight0~56_combout ),
	.datab(portB22),
	.datac(\ShiftRight0~122_combout ),
	.datad(\ShiftRight0~57_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~58 .lut_mask = 16'hFFEA;
defparam \ShiftRight0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N18
cycloneive_lcell_comb \Selector28~5 (
// Equation(s):
// \Selector28~5_combout  = (\Selector3~6_combout  & (!\ShiftRight0~124_combout )) # (!\Selector3~6_combout  & ((\ShiftRight0~124_combout  & (\ShiftRight0~59_combout )) # (!\ShiftRight0~124_combout  & ((\ShiftRight0~58_combout )))))

	.dataa(\Selector3~6_combout ),
	.datab(\ShiftRight0~124_combout ),
	.datac(\ShiftRight0~59_combout ),
	.datad(\ShiftRight0~58_combout ),
	.cin(gnd),
	.combout(\Selector28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~5 .lut_mask = 16'h7362;
defparam \Selector28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N20
cycloneive_lcell_comb \Selector28~6 (
// Equation(s):
// \Selector28~6_combout  = (\Selector3~6_combout  & ((\Selector28~5_combout  & ((\ShiftRight0~64_combout ))) # (!\Selector28~5_combout  & (\ShiftRight0~55_combout )))) # (!\Selector3~6_combout  & (((\Selector28~5_combout ))))

	.dataa(\Selector3~6_combout ),
	.datab(\ShiftRight0~55_combout ),
	.datac(\ShiftRight0~64_combout ),
	.datad(\Selector28~5_combout ),
	.cin(gnd),
	.combout(\Selector28~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~6 .lut_mask = 16'hF588;
defparam \Selector28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N22
cycloneive_lcell_comb \Selector28~8 (
// Equation(s):
// \Selector28~8_combout  = (\Selector28~3_combout ) # ((\Selector28~4_combout ) # ((\Selector28~7_combout  & \Selector28~6_combout )))

	.dataa(\Selector28~3_combout ),
	.datab(\Selector28~7_combout ),
	.datac(\Selector28~4_combout ),
	.datad(\Selector28~6_combout ),
	.cin(gnd),
	.combout(\Selector28~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~8 .lut_mask = 16'hFEFA;
defparam \Selector28~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N10
cycloneive_lcell_comb \ShiftRight0~66 (
// Equation(s):
// \ShiftRight0~66_combout  = (Mux302 & (Mux312 & (\portB~5_combout ))) # (!Mux302 & (!Mux312 & ((\portB~11_combout ))))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB1),
	.datad(portB4),
	.cin(gnd),
	.combout(\ShiftRight0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~66 .lut_mask = 16'h9180;
defparam \ShiftRight0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N0
cycloneive_lcell_comb \ShiftRight0~67 (
// Equation(s):
// \ShiftRight0~67_combout  = (\ShiftRight0~66_combout ) # ((!Mux302 & (Mux312 & \portB~9_combout )))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB3),
	.datad(\ShiftRight0~66_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~67 .lut_mask = 16'hFF40;
defparam \ShiftRight0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N2
cycloneive_lcell_comb \ShiftRight0~68 (
// Equation(s):
// \ShiftRight0~68_combout  = (\ShiftRight0~67_combout ) # ((\portB~7_combout  & \ShiftRight0~122_combout ))

	.dataa(portB2),
	.datab(gnd),
	.datac(\ShiftRight0~122_combout ),
	.datad(\ShiftRight0~67_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~68 .lut_mask = 16'hFFA0;
defparam \ShiftRight0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N0
cycloneive_lcell_comb \ShiftRight0~125 (
// Equation(s):
// \ShiftRight0~125_combout  = (Mux292 & (\ShiftRight0~123_combout  & (\portB~3_combout ))) # (!Mux292 & (((\ShiftRight0~68_combout ))))

	.dataa(\ShiftRight0~123_combout ),
	.datab(Mux292),
	.datac(portB),
	.datad(\ShiftRight0~68_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~125_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~125 .lut_mask = 16'hB380;
defparam \ShiftRight0~125 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N16
cycloneive_lcell_comb \ShiftRight0~72 (
// Equation(s):
// \ShiftRight0~72_combout  = (!Mux302 & ((Mux312 & (\portB~25_combout )) # (!Mux312 & ((\portB~27_combout )))))

	.dataa(Mux302),
	.datab(portB11),
	.datac(Mux312),
	.datad(portB12),
	.cin(gnd),
	.combout(\ShiftRight0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~72 .lut_mask = 16'h4540;
defparam \ShiftRight0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N26
cycloneive_lcell_comb \ShiftRight0~73 (
// Equation(s):
// \ShiftRight0~73_combout  = (Mux302 & ((Mux312 & (\portB~21_combout )) # (!Mux312 & ((\portB~23_combout )))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB9),
	.datad(portB10),
	.cin(gnd),
	.combout(\ShiftRight0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~73 .lut_mask = 16'hC480;
defparam \ShiftRight0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N26
cycloneive_lcell_comb \ShiftRight0~69 (
// Equation(s):
// \ShiftRight0~69_combout  = (!Mux302 & ((Mux312 & ((\portB~17_combout ))) # (!Mux312 & (\portB~19_combout ))))

	.dataa(Mux302),
	.datab(portB8),
	.datac(Mux312),
	.datad(portB7),
	.cin(gnd),
	.combout(\ShiftRight0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~69 .lut_mask = 16'h5404;
defparam \ShiftRight0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N0
cycloneive_lcell_comb \ShiftRight0~70 (
// Equation(s):
// \ShiftRight0~70_combout  = (Mux302 & ((Mux312 & (\portB~13_combout )) # (!Mux312 & ((\portB~15_combout )))))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB5),
	.datad(portB6),
	.cin(gnd),
	.combout(\ShiftRight0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~70 .lut_mask = 16'hA280;
defparam \ShiftRight0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N30
cycloneive_lcell_comb \ShiftRight0~71 (
// Equation(s):
// \ShiftRight0~71_combout  = (\ShiftRight0~69_combout ) # (\ShiftRight0~70_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftRight0~69_combout ),
	.datad(\ShiftRight0~70_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~71 .lut_mask = 16'hFFF0;
defparam \ShiftRight0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N28
cycloneive_lcell_comb \Selector20~0 (
// Equation(s):
// \Selector20~0_combout  = (Mux292 & (((\ShiftRight0~71_combout )))) # (!Mux292 & ((\ShiftRight0~72_combout ) # ((\ShiftRight0~73_combout ))))

	.dataa(Mux292),
	.datab(\ShiftRight0~72_combout ),
	.datac(\ShiftRight0~73_combout ),
	.datad(\ShiftRight0~71_combout ),
	.cin(gnd),
	.combout(\Selector20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~0 .lut_mask = 16'hFE54;
defparam \Selector20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N2
cycloneive_lcell_comb \ShiftRight0~74 (
// Equation(s):
// \ShiftRight0~74_combout  = (Mux28 & (\ShiftRight0~125_combout )) # (!Mux28 & ((\Selector20~0_combout )))

	.dataa(gnd),
	.datab(Mux28),
	.datac(\ShiftRight0~125_combout ),
	.datad(\Selector20~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~74 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N20
cycloneive_lcell_comb \ShiftLeft0~52 (
// Equation(s):
// \ShiftLeft0~52_combout  = (\portB~65_combout  & ((\ShiftRight0~122_combout ) # ((\portB~61_combout  & \ShiftRight0~123_combout )))) # (!\portB~65_combout  & (\portB~61_combout  & (\ShiftRight0~123_combout )))

	.dataa(portB31),
	.datab(portB29),
	.datac(\ShiftRight0~123_combout ),
	.datad(\ShiftRight0~122_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~52 .lut_mask = 16'hEAC0;
defparam \ShiftLeft0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N10
cycloneive_lcell_comb \ShiftLeft0~53 (
// Equation(s):
// \ShiftLeft0~53_combout  = (\ShiftLeft0~52_combout ) # ((Mux312 & (\portB~63_combout  & !Mux302)))

	.dataa(Mux312),
	.datab(portB30),
	.datac(Mux302),
	.datad(\ShiftLeft0~52_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~53 .lut_mask = 16'hFF08;
defparam \ShiftLeft0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N20
cycloneive_lcell_comb \Selector29~0 (
// Equation(s):
// \Selector29~0_combout  = (\portB~61_combout  & ((\Selector0~17_combout ) # ((Mux292 & \Selector0~18_combout ))))

	.dataa(portB29),
	.datab(\Selector0~17_combout ),
	.datac(Mux292),
	.datad(\Selector0~18_combout ),
	.cin(gnd),
	.combout(\Selector29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~0 .lut_mask = 16'hA888;
defparam \Selector29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N14
cycloneive_lcell_comb \Selector29~2 (
// Equation(s):
// \Selector29~2_combout  = (Mux292 & (\Selector0~15_combout  & ((!\portB~61_combout )))) # (!Mux292 & ((\portB~61_combout  & (\Selector0~15_combout )) # (!\portB~61_combout  & ((\Selector0~27_combout )))))

	.dataa(Mux292),
	.datab(\Selector0~15_combout ),
	.datac(\Selector0~27_combout ),
	.datad(portB29),
	.cin(gnd),
	.combout(\Selector29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~2 .lut_mask = 16'h44D8;
defparam \Selector29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N12
cycloneive_lcell_comb \Selector29~1 (
// Equation(s):
// \Selector29~1_combout  = (\Selector0~31_combout  & ((\Add0~4_combout ) # ((\Selector0~14_combout  & \Add1~4_combout )))) # (!\Selector0~31_combout  & (\Selector0~14_combout  & (\Add1~4_combout )))

	.dataa(\Selector0~31_combout ),
	.datab(\Selector0~14_combout ),
	.datac(\Add1~4_combout ),
	.datad(\Add0~4_combout ),
	.cin(gnd),
	.combout(\Selector29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~1 .lut_mask = 16'hEAC0;
defparam \Selector29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N24
cycloneive_lcell_comb \Selector29~3 (
// Equation(s):
// \Selector29~3_combout  = (\Selector29~2_combout ) # ((\Selector29~1_combout ) # ((Mux292 & \Selector0~17_combout )))

	.dataa(Mux292),
	.datab(\Selector29~2_combout ),
	.datac(\Selector0~17_combout ),
	.datad(\Selector29~1_combout ),
	.cin(gnd),
	.combout(\Selector29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~3 .lut_mask = 16'hFFEC;
defparam \Selector29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N30
cycloneive_lcell_comb \ShiftRight0~80 (
// Equation(s):
// \ShiftRight0~80_combout  = (Mux302 & ((Mux312 & ((\portB~39_combout ))) # (!Mux312 & (\portB~41_combout ))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB19),
	.datad(portB18),
	.cin(gnd),
	.combout(\ShiftRight0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~80 .lut_mask = 16'hC840;
defparam \ShiftRight0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N18
cycloneive_lcell_comb \ShiftRight0~77 (
// Equation(s):
// \ShiftRight0~77_combout  = (Mux302 & ((Mux312 & (\portB~31_combout )) # (!Mux312 & ((\portB~33_combout ))))) # (!Mux302 & (((Mux312))))

	.dataa(portB14),
	.datab(portB15),
	.datac(Mux302),
	.datad(Mux312),
	.cin(gnd),
	.combout(\ShiftRight0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~77 .lut_mask = 16'hAFC0;
defparam \ShiftRight0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N28
cycloneive_lcell_comb \ShiftRight0~78 (
// Equation(s):
// \ShiftRight0~78_combout  = (Mux302 & (((\ShiftRight0~77_combout )))) # (!Mux302 & ((\ShiftRight0~77_combout  & ((\portB~35_combout ))) # (!\ShiftRight0~77_combout  & (\portB~37_combout ))))

	.dataa(portB17),
	.datab(Mux302),
	.datac(portB16),
	.datad(\ShiftRight0~77_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~78 .lut_mask = 16'hFC22;
defparam \ShiftRight0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N18
cycloneive_lcell_comb \ShiftRight0~81 (
// Equation(s):
// \ShiftRight0~81_combout  = (Mux292 & (((\ShiftRight0~78_combout )))) # (!Mux292 & ((\ShiftRight0~79_combout ) # ((\ShiftRight0~80_combout ))))

	.dataa(\ShiftRight0~79_combout ),
	.datab(Mux292),
	.datac(\ShiftRight0~80_combout ),
	.datad(\ShiftRight0~78_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~81 .lut_mask = 16'hFE32;
defparam \ShiftRight0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N6
cycloneive_lcell_comb \ShiftRight0~41 (
// Equation(s):
// \ShiftRight0~41_combout  = (Mux312 & (\portB~55_combout )) # (!Mux312 & ((\portB~57_combout )))

	.dataa(gnd),
	.datab(Mux312),
	.datac(portB26),
	.datad(portB27),
	.cin(gnd),
	.combout(\ShiftRight0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~41 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N8
cycloneive_lcell_comb \ShiftRight0~75 (
// Equation(s):
// \ShiftRight0~75_combout  = (Mux312 & (((Mux302 & \portB~47_combout )))) # (!Mux312 & (\portB~53_combout  & (!Mux302)))

	.dataa(portB25),
	.datab(Mux312),
	.datac(Mux302),
	.datad(portB22),
	.cin(gnd),
	.combout(\ShiftRight0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~75 .lut_mask = 16'hC202;
defparam \ShiftRight0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N2
cycloneive_lcell_comb \ShiftRight0~76 (
// Equation(s):
// \ShiftRight0~76_combout  = (\ShiftRight0~75_combout ) # ((\ShiftRight0~52_combout ) # ((\ShiftRight0~122_combout  & \portB~49_combout )))

	.dataa(\ShiftRight0~122_combout ),
	.datab(portB23),
	.datac(\ShiftRight0~75_combout ),
	.datad(\ShiftRight0~52_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~76 .lut_mask = 16'hFFF8;
defparam \ShiftRight0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N24
cycloneive_lcell_comb \Selector29~4 (
// Equation(s):
// \Selector29~4_combout  = (\ShiftRight0~124_combout  & (\ShiftRight0~38_combout  & ((!\Selector3~6_combout )))) # (!\ShiftRight0~124_combout  & (((\ShiftRight0~76_combout ) # (\Selector3~6_combout ))))

	.dataa(\ShiftRight0~38_combout ),
	.datab(\ShiftRight0~124_combout ),
	.datac(\ShiftRight0~76_combout ),
	.datad(\Selector3~6_combout ),
	.cin(gnd),
	.combout(\Selector29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~4 .lut_mask = 16'h33B8;
defparam \Selector29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N12
cycloneive_lcell_comb \Selector29~5 (
// Equation(s):
// \Selector29~5_combout  = (\Selector3~6_combout  & ((\Selector29~4_combout  & (\ShiftRight0~81_combout )) # (!\Selector29~4_combout  & ((\ShiftRight0~41_combout ))))) # (!\Selector3~6_combout  & (((\Selector29~4_combout ))))

	.dataa(\Selector3~6_combout ),
	.datab(\ShiftRight0~81_combout ),
	.datac(\ShiftRight0~41_combout ),
	.datad(\Selector29~4_combout ),
	.cin(gnd),
	.combout(\Selector29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~5 .lut_mask = 16'hDDA0;
defparam \Selector29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N14
cycloneive_lcell_comb \Selector29~6 (
// Equation(s):
// \Selector29~6_combout  = (\Selector29~0_combout ) # ((\Selector29~3_combout ) # ((\Selector28~7_combout  & \Selector29~5_combout )))

	.dataa(\Selector29~0_combout ),
	.datab(\Selector28~7_combout ),
	.datac(\Selector29~3_combout ),
	.datad(\Selector29~5_combout ),
	.cin(gnd),
	.combout(\Selector29~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~6 .lut_mask = 16'hFEFA;
defparam \Selector29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N22
cycloneive_lcell_comb \ShiftRight0~83 (
// Equation(s):
// \ShiftRight0~83_combout  = (Mux302 & (Mux312 & (\portB~7_combout ))) # (!Mux302 & (!Mux312 & ((\portB~13_combout ))))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB2),
	.datad(portB5),
	.cin(gnd),
	.combout(\ShiftRight0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~83 .lut_mask = 16'h9180;
defparam \ShiftRight0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N28
cycloneive_lcell_comb \ShiftRight0~82 (
// Equation(s):
// \ShiftRight0~82_combout  = (Mux312 & (!Mux302 & \portB~11_combout ))

	.dataa(gnd),
	.datab(Mux312),
	.datac(Mux302),
	.datad(portB4),
	.cin(gnd),
	.combout(\ShiftRight0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~82 .lut_mask = 16'h0C00;
defparam \ShiftRight0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N16
cycloneive_lcell_comb \ShiftRight0~84 (
// Equation(s):
// \ShiftRight0~84_combout  = (\ShiftRight0~83_combout ) # ((\ShiftRight0~82_combout ) # ((\portB~9_combout  & \ShiftRight0~122_combout )))

	.dataa(portB3),
	.datab(\ShiftRight0~122_combout ),
	.datac(\ShiftRight0~83_combout ),
	.datad(\ShiftRight0~82_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~84 .lut_mask = 16'hFFF8;
defparam \ShiftRight0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N10
cycloneive_lcell_comb \ShiftRight0~88 (
// Equation(s):
// \ShiftRight0~88_combout  = (!Mux302 & ((Mux312 & ((\portB~27_combout ))) # (!Mux312 & (\portB~29_combout ))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB13),
	.datad(portB12),
	.cin(gnd),
	.combout(\ShiftRight0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~88 .lut_mask = 16'h3210;
defparam \ShiftRight0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N12
cycloneive_lcell_comb \ShiftRight0~86 (
// Equation(s):
// \ShiftRight0~86_combout  = (Mux302 & (\portB~15_combout  & (Mux312))) # (!Mux302 & (((!Mux312 & \portB~21_combout ))))

	.dataa(Mux302),
	.datab(portB6),
	.datac(Mux312),
	.datad(portB9),
	.cin(gnd),
	.combout(\ShiftRight0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~86 .lut_mask = 16'h8580;
defparam \ShiftRight0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N18
cycloneive_lcell_comb \ShiftRight0~87 (
// Equation(s):
// \ShiftRight0~87_combout  = (\ShiftRight0~51_combout ) # ((\ShiftRight0~86_combout ) # ((\ShiftRight0~122_combout  & \portB~17_combout )))

	.dataa(\ShiftRight0~122_combout ),
	.datab(portB7),
	.datac(\ShiftRight0~51_combout ),
	.datad(\ShiftRight0~86_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~87 .lut_mask = 16'hFFF8;
defparam \ShiftRight0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N20
cycloneive_lcell_comb \ShiftRight0~89 (
// Equation(s):
// \ShiftRight0~89_combout  = (Mux302 & ((Mux312 & ((\portB~23_combout ))) # (!Mux312 & (\portB~25_combout ))))

	.dataa(portB11),
	.datab(portB10),
	.datac(Mux302),
	.datad(Mux312),
	.cin(gnd),
	.combout(\ShiftRight0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~89 .lut_mask = 16'hC0A0;
defparam \ShiftRight0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N4
cycloneive_lcell_comb \Selector21~0 (
// Equation(s):
// \Selector21~0_combout  = (Mux292 & (((\ShiftRight0~87_combout )))) # (!Mux292 & ((\ShiftRight0~88_combout ) # ((\ShiftRight0~89_combout ))))

	.dataa(\ShiftRight0~88_combout ),
	.datab(Mux292),
	.datac(\ShiftRight0~87_combout ),
	.datad(\ShiftRight0~89_combout ),
	.cin(gnd),
	.combout(\Selector21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~0 .lut_mask = 16'hF3E2;
defparam \Selector21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N14
cycloneive_lcell_comb \ShiftLeft0~55 (
// Equation(s):
// \ShiftLeft0~55_combout  = (\portB~55_combout  & ((\ShiftRight0~123_combout ) # ((\portB~59_combout  & \ShiftRight0~122_combout )))) # (!\portB~55_combout  & (\portB~59_combout  & ((\ShiftRight0~122_combout ))))

	.dataa(portB26),
	.datab(portB28),
	.datac(\ShiftRight0~123_combout ),
	.datad(\ShiftRight0~122_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~55 .lut_mask = 16'hECA0;
defparam \ShiftLeft0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N24
cycloneive_lcell_comb \ShiftLeft0~54 (
// Equation(s):
// \ShiftLeft0~54_combout  = (Mux312 & ((Mux302 & ((\portB~61_combout ))) # (!Mux302 & (\portB~57_combout ))))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB27),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~54 .lut_mask = 16'hC840;
defparam \ShiftLeft0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N4
cycloneive_lcell_comb \ShiftLeft0~56 (
// Equation(s):
// \ShiftLeft0~56_combout  = (!Mux292 & ((\ShiftLeft0~55_combout ) # (\ShiftLeft0~54_combout )))

	.dataa(Mux292),
	.datab(gnd),
	.datac(\ShiftLeft0~55_combout ),
	.datad(\ShiftLeft0~54_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~56 .lut_mask = 16'h5550;
defparam \ShiftLeft0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N22
cycloneive_lcell_comb \ShiftLeft0~61 (
// Equation(s):
// \ShiftLeft0~61_combout  = (\portB~43_combout  & ((\ShiftRight0~122_combout ) # ((\ShiftRight0~123_combout  & \portB~39_combout )))) # (!\portB~43_combout  & (((\ShiftRight0~123_combout  & \portB~39_combout ))))

	.dataa(portB20),
	.datab(\ShiftRight0~122_combout ),
	.datac(\ShiftRight0~123_combout ),
	.datad(portB18),
	.cin(gnd),
	.combout(\ShiftLeft0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~61 .lut_mask = 16'hF888;
defparam \ShiftLeft0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N16
cycloneive_lcell_comb \ShiftLeft0~58 (
// Equation(s):
// \ShiftLeft0~58_combout  = (Mux302 & ((Mux312 & (\portB~53_combout )) # (!Mux312 & ((\portB~51_combout )))))

	.dataa(portB25),
	.datab(Mux312),
	.datac(Mux302),
	.datad(portB24),
	.cin(gnd),
	.combout(\ShiftLeft0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~58 .lut_mask = 16'hB080;
defparam \ShiftLeft0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N14
cycloneive_lcell_comb \ShiftLeft0~59 (
// Equation(s):
// \ShiftLeft0~59_combout  = (\ShiftRight0~56_combout ) # ((\ShiftLeft0~58_combout ) # ((\ShiftRight0~123_combout  & \portB~47_combout )))

	.dataa(\ShiftRight0~56_combout ),
	.datab(\ShiftRight0~123_combout ),
	.datac(portB22),
	.datad(\ShiftLeft0~58_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~59 .lut_mask = 16'hFFEA;
defparam \ShiftLeft0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N14
cycloneive_lcell_comb \ShiftLeft0~60 (
// Equation(s):
// \ShiftLeft0~60_combout  = (Mux312 & ((Mux302 & (\portB~45_combout )) # (!Mux302 & ((\portB~41_combout )))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB21),
	.datad(portB19),
	.cin(gnd),
	.combout(\ShiftLeft0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~60 .lut_mask = 16'hA280;
defparam \ShiftLeft0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N24
cycloneive_lcell_comb \Selector10~0 (
// Equation(s):
// \Selector10~0_combout  = (Mux292 & (((\ShiftLeft0~59_combout )))) # (!Mux292 & ((\ShiftLeft0~61_combout ) # ((\ShiftLeft0~60_combout ))))

	.dataa(\ShiftLeft0~61_combout ),
	.datab(Mux292),
	.datac(\ShiftLeft0~59_combout ),
	.datad(\ShiftLeft0~60_combout ),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~0 .lut_mask = 16'hF3E2;
defparam \Selector10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N8
cycloneive_lcell_comb \Selector10~2 (
// Equation(s):
// \Selector10~2_combout  = (\Selector0~14_combout  & ((\Add1~42_combout ) # ((\Selector0~31_combout  & \Add0~42_combout )))) # (!\Selector0~14_combout  & (\Selector0~31_combout  & ((\Add0~42_combout ))))

	.dataa(\Selector0~14_combout ),
	.datab(\Selector0~31_combout ),
	.datac(\Add1~42_combout ),
	.datad(\Add0~42_combout ),
	.cin(gnd),
	.combout(\Selector10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~2 .lut_mask = 16'hECA0;
defparam \Selector10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N0
cycloneive_lcell_comb \Selector10~3 (
// Equation(s):
// \Selector10~3_combout  = (\portB~23_combout  & ((\Selector0~17_combout ) # ((Mux10 & \Selector0~18_combout ))))

	.dataa(Mux10),
	.datab(\Selector0~17_combout ),
	.datac(portB10),
	.datad(\Selector0~18_combout ),
	.cin(gnd),
	.combout(\Selector10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~3 .lut_mask = 16'hE0C0;
defparam \Selector10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N22
cycloneive_lcell_comb \Selector10~4 (
// Equation(s):
// \Selector10~4_combout  = (\Selector10~3_combout ) # ((!Mux10 & (\Selector0~27_combout  & !\portB~23_combout )))

	.dataa(Mux10),
	.datab(\Selector0~27_combout ),
	.datac(portB10),
	.datad(\Selector10~3_combout ),
	.cin(gnd),
	.combout(\Selector10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~4 .lut_mask = 16'hFF04;
defparam \Selector10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N22
cycloneive_lcell_comb \Selector10~5 (
// Equation(s):
// \Selector10~5_combout  = (\Selector10~4_combout ) # ((\Selector0~15_combout  & (Mux10 $ (\portB~23_combout ))))

	.dataa(Mux10),
	.datab(portB10),
	.datac(\Selector10~4_combout ),
	.datad(\Selector0~15_combout ),
	.cin(gnd),
	.combout(\Selector10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~5 .lut_mask = 16'hF6F0;
defparam \Selector10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N0
cycloneive_lcell_comb \ShiftRight0~97 (
// Equation(s):
// \ShiftRight0~97_combout  = (!Mux302 & ((Mux312 & ((\portB~5_combout ))) # (!Mux312 & (\portB~7_combout ))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB2),
	.datad(portB1),
	.cin(gnd),
	.combout(\ShiftRight0~97_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~97 .lut_mask = 16'h3210;
defparam \ShiftRight0~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N30
cycloneive_lcell_comb \ShiftRight0~98 (
// Equation(s):
// \ShiftRight0~98_combout  = (\ShiftRight0~97_combout ) # ((\ShiftRight0~122_combout  & \portB~3_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~122_combout ),
	.datac(portB),
	.datad(\ShiftRight0~97_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~98_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~98 .lut_mask = 16'hFFC0;
defparam \ShiftRight0~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N20
cycloneive_lcell_comb \ShiftRight0~94 (
// Equation(s):
// \ShiftRight0~94_combout  = (Mux302 & ((Mux312 & (\portB~17_combout )) # (!Mux312 & ((\portB~19_combout ))))) # (!Mux302 & (((Mux312))))

	.dataa(Mux302),
	.datab(portB7),
	.datac(Mux312),
	.datad(portB8),
	.cin(gnd),
	.combout(\ShiftRight0~94_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~94 .lut_mask = 16'hDAD0;
defparam \ShiftRight0~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N6
cycloneive_lcell_comb \ShiftRight0~95 (
// Equation(s):
// \ShiftRight0~95_combout  = (Mux302 & (((\ShiftRight0~94_combout )))) # (!Mux302 & ((\ShiftRight0~94_combout  & (\portB~21_combout )) # (!\ShiftRight0~94_combout  & ((\portB~23_combout )))))

	.dataa(Mux302),
	.datab(portB9),
	.datac(portB10),
	.datad(\ShiftRight0~94_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~95_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~95 .lut_mask = 16'hEE50;
defparam \ShiftRight0~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N14
cycloneive_lcell_comb \ShiftRight0~96 (
// Equation(s):
// \ShiftRight0~96_combout  = (\ShiftRight0~93_combout  & ((\Selector7~19_combout ) # ((\ShiftRight0~124_combout  & \ShiftRight0~95_combout )))) # (!\ShiftRight0~93_combout  & (\ShiftRight0~124_combout  & ((\ShiftRight0~95_combout ))))

	.dataa(\ShiftRight0~93_combout ),
	.datab(\ShiftRight0~124_combout ),
	.datac(\Selector7~19_combout ),
	.datad(\ShiftRight0~95_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~96_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~96 .lut_mask = 16'hECA0;
defparam \ShiftRight0~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N14
cycloneive_lcell_comb \ShiftRight0~99 (
// Equation(s):
// \ShiftRight0~99_combout  = (\ShiftRight0~96_combout ) # ((!Mux292 & (Mux28 & \ShiftRight0~98_combout )))

	.dataa(Mux292),
	.datab(Mux28),
	.datac(\ShiftRight0~98_combout ),
	.datad(\ShiftRight0~96_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~99_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~99 .lut_mask = 16'hFF40;
defparam \ShiftRight0~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N30
cycloneive_lcell_comb \ShiftLeft0~63 (
// Equation(s):
// \ShiftLeft0~63_combout  = (\portB~35_combout  & ((\ShiftRight0~122_combout ) # ((\ShiftRight0~123_combout  & \portB~31_combout )))) # (!\portB~35_combout  & (\ShiftRight0~123_combout  & ((\portB~31_combout ))))

	.dataa(portB16),
	.datab(\ShiftRight0~123_combout ),
	.datac(\ShiftRight0~122_combout ),
	.datad(portB14),
	.cin(gnd),
	.combout(\ShiftLeft0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~63 .lut_mask = 16'hECA0;
defparam \ShiftLeft0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N26
cycloneive_lcell_comb \ShiftLeft0~66 (
// Equation(s):
// \ShiftLeft0~66_combout  = (\portB~23_combout  & ((\ShiftRight0~123_combout ) # ((\ShiftRight0~122_combout  & \portB~27_combout )))) # (!\portB~23_combout  & (((\ShiftRight0~122_combout  & \portB~27_combout ))))

	.dataa(portB10),
	.datab(\ShiftRight0~123_combout ),
	.datac(\ShiftRight0~122_combout ),
	.datad(portB12),
	.cin(gnd),
	.combout(\ShiftLeft0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~66 .lut_mask = 16'hF888;
defparam \ShiftLeft0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N28
cycloneive_lcell_comb \ShiftLeft0~65 (
// Equation(s):
// \ShiftLeft0~65_combout  = (Mux312 & ((Mux302 & (\portB~29_combout )) # (!Mux302 & ((\portB~25_combout )))))

	.dataa(portB13),
	.datab(Mux312),
	.datac(Mux302),
	.datad(portB11),
	.cin(gnd),
	.combout(\ShiftLeft0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~65 .lut_mask = 16'h8C80;
defparam \ShiftLeft0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N8
cycloneive_lcell_comb \ShiftLeft0~67 (
// Equation(s):
// \ShiftLeft0~67_combout  = (\ShiftLeft0~66_combout ) # (\ShiftLeft0~65_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftLeft0~66_combout ),
	.datad(\ShiftLeft0~65_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~67 .lut_mask = 16'hFFF0;
defparam \ShiftLeft0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N16
cycloneive_lcell_comb \ShiftLeft0~62 (
// Equation(s):
// \ShiftLeft0~62_combout  = (Mux312 & ((Mux302 & ((\portB~37_combout ))) # (!Mux302 & (\portB~33_combout ))))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB15),
	.datad(portB17),
	.cin(gnd),
	.combout(\ShiftLeft0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~62 .lut_mask = 16'hC840;
defparam \ShiftLeft0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N2
cycloneive_lcell_comb \ShiftLeft0~103 (
// Equation(s):
// \ShiftLeft0~103_combout  = (Mux292 & ((\ShiftLeft0~63_combout ) # ((\ShiftLeft0~62_combout )))) # (!Mux292 & (((\ShiftLeft0~67_combout ))))

	.dataa(\ShiftLeft0~63_combout ),
	.datab(Mux292),
	.datac(\ShiftLeft0~67_combout ),
	.datad(\ShiftLeft0~62_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~103_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~103 .lut_mask = 16'hFCB8;
defparam \ShiftLeft0~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N28
cycloneive_lcell_comb \Selector2~7 (
// Equation(s):
// \Selector2~7_combout  = (\portB~7_combout  & (\Selector0~15_combout  & ((!Mux2)))) # (!\portB~7_combout  & ((Mux2 & (\Selector0~15_combout )) # (!Mux2 & ((\Selector0~27_combout )))))

	.dataa(\Selector0~15_combout ),
	.datab(portB2),
	.datac(\Selector0~27_combout ),
	.datad(Mux2),
	.cin(gnd),
	.combout(\Selector2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~7 .lut_mask = 16'h22B8;
defparam \Selector2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N26
cycloneive_lcell_comb \Selector2~8 (
// Equation(s):
// \Selector2~8_combout  = (\Selector2~7_combout ) # ((\ShiftRight0~124_combout  & (\ShiftRight0~98_combout  & Selector8)))

	.dataa(\ShiftRight0~124_combout ),
	.datab(\Selector2~7_combout ),
	.datac(\ShiftRight0~98_combout ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Selector2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~8 .lut_mask = 16'hECCC;
defparam \Selector2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N22
cycloneive_lcell_comb \ShiftLeft0~68 (
// Equation(s):
// \ShiftLeft0~68_combout  = (Mux312 & ((Mux302 & ((\portB~21_combout ))) # (!Mux302 & (\portB~17_combout ))))

	.dataa(Mux302),
	.datab(portB7),
	.datac(Mux312),
	.datad(portB9),
	.cin(gnd),
	.combout(\ShiftLeft0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~68 .lut_mask = 16'hE040;
defparam \ShiftLeft0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N12
cycloneive_lcell_comb \ShiftLeft0~69 (
// Equation(s):
// \ShiftLeft0~69_combout  = (\ShiftRight0~122_combout  & ((\portB~19_combout ) # ((\ShiftRight0~123_combout  & \portB~15_combout )))) # (!\ShiftRight0~122_combout  & (\ShiftRight0~123_combout  & (\portB~15_combout )))

	.dataa(\ShiftRight0~122_combout ),
	.datab(\ShiftRight0~123_combout ),
	.datac(portB6),
	.datad(portB8),
	.cin(gnd),
	.combout(\ShiftLeft0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~69 .lut_mask = 16'hEAC0;
defparam \ShiftLeft0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N10
cycloneive_lcell_comb \ShiftLeft0~70 (
// Equation(s):
// \ShiftLeft0~70_combout  = (\ShiftLeft0~68_combout ) # (\ShiftLeft0~69_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftLeft0~68_combout ),
	.datad(\ShiftLeft0~69_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~70 .lut_mask = 16'hFFF0;
defparam \ShiftLeft0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N0
cycloneive_lcell_comb \Selector2~1 (
// Equation(s):
// \Selector2~1_combout  = (\ShiftRight0~124_combout  & (\ShiftLeft0~14_combout  & (!\Selector3~6_combout ))) # (!\ShiftRight0~124_combout  & (((\Selector3~6_combout ) # (\ShiftLeft0~70_combout ))))

	.dataa(\ShiftLeft0~14_combout ),
	.datab(\ShiftRight0~124_combout ),
	.datac(\Selector3~6_combout ),
	.datad(\ShiftLeft0~70_combout ),
	.cin(gnd),
	.combout(\Selector2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~1 .lut_mask = 16'h3B38;
defparam \Selector2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N18
cycloneive_lcell_comb \Selector2~2 (
// Equation(s):
// \Selector2~2_combout  = (\Selector2~1_combout  & (((\ShiftLeft0~103_combout ) # (!\Selector3~6_combout )))) # (!\Selector2~1_combout  & (\ShiftLeft0~16_combout  & (\Selector3~6_combout )))

	.dataa(\ShiftLeft0~16_combout ),
	.datab(\Selector2~1_combout ),
	.datac(\Selector3~6_combout ),
	.datad(\ShiftLeft0~103_combout ),
	.cin(gnd),
	.combout(\Selector2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~2 .lut_mask = 16'hEC2C;
defparam \Selector2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N20
cycloneive_lcell_comb \Selector2~5 (
// Equation(s):
// \Selector2~5_combout  = (\Selector0~17_combout  & (((Mux2) # (\portB~7_combout )))) # (!\Selector0~17_combout  & (\Selector0~18_combout  & (Mux2 & \portB~7_combout )))

	.dataa(\Selector0~17_combout ),
	.datab(\Selector0~18_combout ),
	.datac(Mux2),
	.datad(portB2),
	.cin(gnd),
	.combout(\Selector2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~5 .lut_mask = 16'hEAA0;
defparam \Selector2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N26
cycloneive_lcell_comb \Selector2~3 (
// Equation(s):
// \Selector2~3_combout  = (\Selector1~11_combout  & ((Mux28 & (ShiftLeft0)) # (!Mux28 & ((\Selector10~0_combout )))))

	.dataa(Mux28),
	.datab(ShiftLeft0),
	.datac(\Selector10~0_combout ),
	.datad(\Selector1~11_combout ),
	.cin(gnd),
	.combout(\Selector2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~3 .lut_mask = 16'hD800;
defparam \Selector2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N4
cycloneive_lcell_comb \Selector2~4 (
// Equation(s):
// \Selector2~4_combout  = (\Selector2~3_combout ) # ((\Selector0~31_combout  & \Add0~58_combout ))

	.dataa(\Selector0~31_combout ),
	.datab(gnd),
	.datac(\Selector2~3_combout ),
	.datad(\Add0~58_combout ),
	.cin(gnd),
	.combout(\Selector2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~4 .lut_mask = 16'hFAF0;
defparam \Selector2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N2
cycloneive_lcell_comb \Selector2~6 (
// Equation(s):
// \Selector2~6_combout  = (\Selector2~5_combout ) # ((\Selector2~4_combout ) # ((\Selector2~2_combout  & \Selector2~0_combout )))

	.dataa(\Selector2~2_combout ),
	.datab(\Selector2~5_combout ),
	.datac(\Selector2~4_combout ),
	.datad(\Selector2~0_combout ),
	.cin(gnd),
	.combout(\Selector2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~6 .lut_mask = 16'hFEFC;
defparam \Selector2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N14
cycloneive_lcell_comb \Selector1~16 (
// Equation(s):
// \Selector1~16_combout  = (!Mux1 & (\Selector0~27_combout  & !\portB~5_combout ))

	.dataa(gnd),
	.datab(Mux1),
	.datac(\Selector0~27_combout ),
	.datad(portB1),
	.cin(gnd),
	.combout(\Selector1~16_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~16 .lut_mask = 16'h0030;
defparam \Selector1~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N16
cycloneive_lcell_comb \Selector1~17 (
// Equation(s):
// \Selector1~17_combout  = (\Selector1~26_combout  & ((\Selector0~22_combout ) # ((Mux1 & \Selector0~17_combout )))) # (!\Selector1~26_combout  & (Mux1 & (\Selector0~17_combout )))

	.dataa(\Selector1~26_combout ),
	.datab(Mux1),
	.datac(\Selector0~17_combout ),
	.datad(\Selector0~22_combout ),
	.cin(gnd),
	.combout(\Selector1~17_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~17 .lut_mask = 16'hEAC0;
defparam \Selector1~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N26
cycloneive_lcell_comb \Selector1~18 (
// Equation(s):
// \Selector1~18_combout  = (\Selector1~16_combout ) # ((\Selector1~17_combout ) # ((\Selector0~31_combout  & \Add0~60_combout )))

	.dataa(\Selector0~31_combout ),
	.datab(\Selector1~16_combout ),
	.datac(\Add0~60_combout ),
	.datad(\Selector1~17_combout ),
	.cin(gnd),
	.combout(\Selector1~18_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~18 .lut_mask = 16'hFFEC;
defparam \Selector1~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N20
cycloneive_lcell_comb \ShiftLeft0~71 (
// Equation(s):
// \ShiftLeft0~71_combout  = (Mux312 & (!Mux302 & \portB~55_combout ))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(gnd),
	.datad(portB26),
	.cin(gnd),
	.combout(\ShiftLeft0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~71 .lut_mask = 16'h2200;
defparam \ShiftLeft0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N6
cycloneive_lcell_comb \ShiftLeft0~72 (
// Equation(s):
// \ShiftLeft0~72_combout  = (Mux302 & ((Mux312 & ((\portB~59_combout ))) # (!Mux312 & (\portB~57_combout ))))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB27),
	.datad(portB28),
	.cin(gnd),
	.combout(\ShiftLeft0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~72 .lut_mask = 16'hA820;
defparam \ShiftLeft0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N14
cycloneive_lcell_comb \ShiftLeft0~73 (
// Equation(s):
// \ShiftLeft0~73_combout  = (\ShiftLeft0~71_combout ) # ((\ShiftLeft0~72_combout ) # ((\portB~53_combout  & \ShiftRight0~123_combout )))

	.dataa(portB25),
	.datab(\ShiftLeft0~71_combout ),
	.datac(\ShiftRight0~123_combout ),
	.datad(\ShiftLeft0~72_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~73 .lut_mask = 16'hFFEC;
defparam \ShiftLeft0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N8
cycloneive_lcell_comb \ShiftLeft0~74 (
// Equation(s):
// \ShiftLeft0~74_combout  = (Mux292 & ((\ShiftLeft0~53_combout ))) # (!Mux292 & (\ShiftLeft0~73_combout ))

	.dataa(Mux292),
	.datab(gnd),
	.datac(\ShiftLeft0~73_combout ),
	.datad(\ShiftLeft0~53_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~74 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N10
cycloneive_lcell_comb \ShiftLeft0~75 (
// Equation(s):
// \ShiftLeft0~75_combout  = (Mux312 & ((Mux302 & ((\portB~51_combout ))) # (!Mux302 & (\portB~47_combout ))))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB22),
	.datad(portB24),
	.cin(gnd),
	.combout(\ShiftLeft0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~75 .lut_mask = 16'hC840;
defparam \ShiftLeft0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N10
cycloneive_lcell_comb \ShiftLeft0~76 (
// Equation(s):
// \ShiftLeft0~76_combout  = (\portB~45_combout  & ((\ShiftRight0~123_combout ) # ((\ShiftRight0~122_combout  & \portB~49_combout )))) # (!\portB~45_combout  & (\ShiftRight0~122_combout  & ((\portB~49_combout ))))

	.dataa(portB21),
	.datab(\ShiftRight0~122_combout ),
	.datac(\ShiftRight0~123_combout ),
	.datad(portB23),
	.cin(gnd),
	.combout(\ShiftLeft0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~76 .lut_mask = 16'hECA0;
defparam \ShiftLeft0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N4
cycloneive_lcell_comb \ShiftLeft0~77 (
// Equation(s):
// \ShiftLeft0~77_combout  = (\ShiftLeft0~75_combout ) # (\ShiftLeft0~76_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftLeft0~75_combout ),
	.datad(\ShiftLeft0~76_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~77 .lut_mask = 16'hFFF0;
defparam \ShiftLeft0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N30
cycloneive_lcell_comb \ShiftLeft0~79 (
// Equation(s):
// \ShiftLeft0~79_combout  = (\portB~37_combout  & ((\ShiftRight0~123_combout ) # ((\ShiftRight0~122_combout  & \portB~41_combout )))) # (!\portB~37_combout  & (\ShiftRight0~122_combout  & ((\portB~41_combout ))))

	.dataa(portB17),
	.datab(\ShiftRight0~122_combout ),
	.datac(\ShiftRight0~123_combout ),
	.datad(portB19),
	.cin(gnd),
	.combout(\ShiftLeft0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~79 .lut_mask = 16'hECA0;
defparam \ShiftLeft0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N30
cycloneive_lcell_comb \ShiftLeft0~78 (
// Equation(s):
// \ShiftLeft0~78_combout  = (Mux312 & ((Mux302 & (\portB~43_combout )) # (!Mux302 & ((\portB~39_combout )))))

	.dataa(portB20),
	.datab(Mux312),
	.datac(Mux302),
	.datad(portB18),
	.cin(gnd),
	.combout(\ShiftLeft0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~78 .lut_mask = 16'h8C80;
defparam \ShiftLeft0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N28
cycloneive_lcell_comb \Selector9~0 (
// Equation(s):
// \Selector9~0_combout  = (Mux292 & (\ShiftLeft0~77_combout )) # (!Mux292 & (((\ShiftLeft0~79_combout ) # (\ShiftLeft0~78_combout ))))

	.dataa(Mux292),
	.datab(\ShiftLeft0~77_combout ),
	.datac(\ShiftLeft0~79_combout ),
	.datad(\ShiftLeft0~78_combout ),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~0 .lut_mask = 16'hDDD8;
defparam \Selector9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N18
cycloneive_lcell_comb \Selector1~12 (
// Equation(s):
// \Selector1~12_combout  = (\Selector1~11_combout  & ((Mux28 & (\ShiftLeft0~74_combout )) # (!Mux28 & ((\Selector9~0_combout )))))

	.dataa(\ShiftLeft0~74_combout ),
	.datab(Mux28),
	.datac(\Selector9~0_combout ),
	.datad(\Selector1~11_combout ),
	.cin(gnd),
	.combout(\Selector1~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~12 .lut_mask = 16'hB800;
defparam \Selector1~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N28
cycloneive_lcell_comb \Selector1~22 (
// Equation(s):
// \Selector1~22_combout  = (\Selector0~15_combout  & (\portB~5_combout  $ (Mux1)))

	.dataa(portB1),
	.datab(Mux1),
	.datac(gnd),
	.datad(\Selector0~15_combout ),
	.cin(gnd),
	.combout(\Selector1~22_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~22 .lut_mask = 16'h6600;
defparam \Selector1~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N12
cycloneive_lcell_comb \Selector1~20 (
// Equation(s):
// \Selector1~20_combout  = (!Mux292 & (!Mux28 & !Mux302))

	.dataa(Mux292),
	.datab(Mux28),
	.datac(gnd),
	.datad(Mux302),
	.cin(gnd),
	.combout(\Selector1~20_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~20 .lut_mask = 16'h0011;
defparam \Selector1~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N8
cycloneive_lcell_comb \Selector1~19 (
// Equation(s):
// \Selector1~19_combout  = (\portB~5_combout  & ((\Selector0~17_combout ) # ((Mux1 & \Selector0~18_combout ))))

	.dataa(\Selector0~17_combout ),
	.datab(Mux1),
	.datac(\Selector0~18_combout ),
	.datad(portB1),
	.cin(gnd),
	.combout(\Selector1~19_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~19 .lut_mask = 16'hEA00;
defparam \Selector1~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N18
cycloneive_lcell_comb \Selector1~21 (
// Equation(s):
// \Selector1~21_combout  = (\Selector1~19_combout ) # ((\ShiftRight0~25_combout  & (\Selector1~20_combout  & Selector8)))

	.dataa(\ShiftRight0~25_combout ),
	.datab(\Selector1~20_combout ),
	.datac(\Selector1~19_combout ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Selector1~21_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~21 .lut_mask = 16'hF8F0;
defparam \Selector1~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N2
cycloneive_lcell_comb \Selector1~23 (
// Equation(s):
// \Selector1~23_combout  = (\Selector1~22_combout ) # ((\Selector1~21_combout ) # ((\Selector0~14_combout  & \Add1~60_combout )))

	.dataa(\Selector0~14_combout ),
	.datab(\Selector1~22_combout ),
	.datac(\Add1~60_combout ),
	.datad(\Selector1~21_combout ),
	.cin(gnd),
	.combout(\Selector1~23_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~23 .lut_mask = 16'hFFEC;
defparam \Selector1~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N30
cycloneive_lcell_comb \ShiftLeft0~32 (
// Equation(s):
// \ShiftLeft0~32_combout  = (Mux312 & ((\portB~11_combout ))) # (!Mux312 & (\portB~9_combout ))

	.dataa(gnd),
	.datab(Mux312),
	.datac(portB3),
	.datad(portB4),
	.cin(gnd),
	.combout(\ShiftLeft0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~32 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N8
cycloneive_lcell_comb \Selector1~13 (
// Equation(s):
// \Selector1~13_combout  = (\Selector1~25_combout  & ((\Selector1~10_combout ) # ((\ShiftLeft0~32_combout )))) # (!\Selector1~25_combout  & (!\Selector1~10_combout  & (\portB~5_combout )))

	.dataa(\Selector1~25_combout ),
	.datab(\Selector1~10_combout ),
	.datac(portB1),
	.datad(\ShiftLeft0~32_combout ),
	.cin(gnd),
	.combout(\Selector1~13_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~13 .lut_mask = 16'hBA98;
defparam \Selector1~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N10
cycloneive_lcell_comb \ShiftLeft0~80 (
// Equation(s):
// \ShiftLeft0~80_combout  = (Mux302 & ((Mux312 & ((\portB~19_combout ))) # (!Mux312 & (\portB~17_combout ))))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB7),
	.datad(portB8),
	.cin(gnd),
	.combout(\ShiftLeft0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~80 .lut_mask = 16'hA820;
defparam \ShiftLeft0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N30
cycloneive_lcell_comb \ShiftLeft0~81 (
// Equation(s):
// \ShiftLeft0~81_combout  = (\ShiftLeft0~80_combout ) # ((!Mux302 & \ShiftLeft0~29_combout ))

	.dataa(Mux302),
	.datab(gnd),
	.datac(\ShiftLeft0~80_combout ),
	.datad(\ShiftLeft0~29_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~81 .lut_mask = 16'hF5F0;
defparam \ShiftLeft0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N18
cycloneive_lcell_comb \Selector1~14 (
// Equation(s):
// \Selector1~14_combout  = (\Selector1~10_combout  & ((\Selector1~13_combout  & ((\ShiftLeft0~81_combout ))) # (!\Selector1~13_combout  & (\portB~7_combout )))) # (!\Selector1~10_combout  & (((\Selector1~13_combout ))))

	.dataa(portB2),
	.datab(\Selector1~10_combout ),
	.datac(\Selector1~13_combout ),
	.datad(\ShiftLeft0~81_combout ),
	.cin(gnd),
	.combout(\Selector1~14_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~14 .lut_mask = 16'hF838;
defparam \Selector1~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N20
cycloneive_lcell_comb \Selector1~15 (
// Equation(s):
// \Selector1~15_combout  = (\Selector16~0_combout  & (!cuifALUOP_0 & \Selector1~14_combout ))

	.dataa(gnd),
	.datab(\Selector16~0_combout ),
	.datac(cuifALUOP_0),
	.datad(\Selector1~14_combout ),
	.cin(gnd),
	.combout(\Selector1~15_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~15 .lut_mask = 16'h0C00;
defparam \Selector1~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N10
cycloneive_lcell_comb \Selector0~7 (
// Equation(s):
// \Selector0~7_combout  = (cuifALUOP_1 & (cuifALUOP_0 & (!cuifALUOP_3 & cuifALUOP_2)))

	.dataa(cuifALUOP_1),
	.datab(cuifALUOP_0),
	.datac(cuifALUOP_3),
	.datad(cuifALUOP_2),
	.cin(gnd),
	.combout(\Selector0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~7 .lut_mask = 16'h0800;
defparam \Selector0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N6
cycloneive_lcell_comb \Selector4~7 (
// Equation(s):
// \Selector4~7_combout  = (\portB~11_combout  & ((\Selector0~5_combout ) # ((Mux4 & \Selector0~6_combout ))))

	.dataa(Mux4),
	.datab(\Selector0~5_combout ),
	.datac(portB4),
	.datad(\Selector0~6_combout ),
	.cin(gnd),
	.combout(\Selector4~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~7 .lut_mask = 16'hE0C0;
defparam \Selector4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N28
cycloneive_lcell_comb \Selector4~8 (
// Equation(s):
// \Selector4~8_combout  = (\Selector4~7_combout ) # ((!\portB~11_combout  & (\Selector0~7_combout  & !Mux4)))

	.dataa(portB4),
	.datab(\Selector0~7_combout ),
	.datac(Mux4),
	.datad(\Selector4~7_combout ),
	.cin(gnd),
	.combout(\Selector4~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~8 .lut_mask = 16'hFF04;
defparam \Selector4~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N2
cycloneive_lcell_comb \Selector4~9 (
// Equation(s):
// \Selector4~9_combout  = (\Selector4~8_combout ) # ((\Selector0~11_combout  & (Mux4 $ (\portB~11_combout ))))

	.dataa(Mux4),
	.datab(\Selector0~11_combout ),
	.datac(portB4),
	.datad(\Selector4~8_combout ),
	.cin(gnd),
	.combout(\Selector4~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~9 .lut_mask = 16'hFF48;
defparam \Selector4~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N2
cycloneive_lcell_comb \ShiftLeft0~24 (
// Equation(s):
// \ShiftLeft0~24_combout  = (Mux312 & ((Mux302 & (\portB~49_combout )) # (!Mux302 & ((\portB~45_combout )))))

	.dataa(Mux312),
	.datab(portB23),
	.datac(portB21),
	.datad(Mux302),
	.cin(gnd),
	.combout(\ShiftLeft0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~24 .lut_mask = 16'h88A0;
defparam \ShiftLeft0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N24
cycloneive_lcell_comb \ShiftLeft0~26 (
// Equation(s):
// \ShiftLeft0~26_combout  = (\ShiftLeft0~25_combout ) # (\ShiftLeft0~24_combout )

	.dataa(\ShiftLeft0~25_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ShiftLeft0~24_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~26 .lut_mask = 16'hFFAA;
defparam \ShiftLeft0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N28
cycloneive_lcell_comb \ShiftLeft0~89 (
// Equation(s):
// \ShiftLeft0~89_combout  = (\ShiftLeft0~23_combout  & ((\Selector7~19_combout ) # ((\ShiftRight0~124_combout  & \ShiftLeft0~26_combout )))) # (!\ShiftLeft0~23_combout  & (\ShiftRight0~124_combout  & ((\ShiftLeft0~26_combout ))))

	.dataa(\ShiftLeft0~23_combout ),
	.datab(\ShiftRight0~124_combout ),
	.datac(\Selector7~19_combout ),
	.datad(\ShiftLeft0~26_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~89 .lut_mask = 16'hECA0;
defparam \ShiftLeft0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N6
cycloneive_lcell_comb \ShiftLeft0~90 (
// Equation(s):
// \ShiftLeft0~90_combout  = (\ShiftLeft0~89_combout ) # ((\ShiftLeft0~20_combout  & (!Mux292 & Mux28)))

	.dataa(\ShiftLeft0~20_combout ),
	.datab(Mux292),
	.datac(Mux28),
	.datad(\ShiftLeft0~89_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~90_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~90 .lut_mask = 16'hFF20;
defparam \ShiftLeft0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N12
cycloneive_lcell_comb \Selector4~4 (
// Equation(s):
// \Selector4~4_combout  = (\Selector7~10_combout  & ((\Selector7~18_combout ) # ((\ShiftLeft0~13_combout )))) # (!\Selector7~10_combout  & (!\Selector7~18_combout  & ((\ShiftLeft0~17_combout ))))

	.dataa(\Selector7~10_combout ),
	.datab(\Selector7~18_combout ),
	.datac(\ShiftLeft0~13_combout ),
	.datad(\ShiftLeft0~17_combout ),
	.cin(gnd),
	.combout(\Selector4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~4 .lut_mask = 16'hB9A8;
defparam \Selector4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N30
cycloneive_lcell_comb \Selector4~5 (
// Equation(s):
// \Selector4~5_combout  = (\Selector7~18_combout  & ((\Selector4~4_combout  & ((\ShiftLeft0~90_combout ))) # (!\Selector4~4_combout  & (\ShiftLeft0~88_combout )))) # (!\Selector7~18_combout  & (((\Selector4~4_combout ))))

	.dataa(\ShiftLeft0~88_combout ),
	.datab(\Selector7~18_combout ),
	.datac(\ShiftLeft0~90_combout ),
	.datad(\Selector4~4_combout ),
	.cin(gnd),
	.combout(\Selector4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~5 .lut_mask = 16'hF388;
defparam \Selector4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N6
cycloneive_lcell_comb \Selector4~2 (
// Equation(s):
// \Selector4~2_combout  = (\Selector0~10_combout  & ((\Add0~54_combout ) # ((\Selector0~8_combout  & \Add1~54_combout )))) # (!\Selector0~10_combout  & (\Selector0~8_combout  & (\Add1~54_combout )))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~8_combout ),
	.datac(\Add1~54_combout ),
	.datad(\Add0~54_combout ),
	.cin(gnd),
	.combout(\Selector4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~2 .lut_mask = 16'hEAC0;
defparam \Selector4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N12
cycloneive_lcell_comb \Selector4~3 (
// Equation(s):
// \Selector4~3_combout  = (\Selector4~2_combout ) # ((Mux4 & \Selector0~5_combout ))

	.dataa(Mux4),
	.datab(gnd),
	.datac(\Selector0~5_combout ),
	.datad(\Selector4~2_combout ),
	.cin(gnd),
	.combout(\Selector4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~3 .lut_mask = 16'hFFA0;
defparam \Selector4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N16
cycloneive_lcell_comb \Selector4~6 (
// Equation(s):
// \Selector4~6_combout  = (\Selector4~3_combout ) # ((!\ShiftRight0~22_combout  & (\Selector0~9_combout  & \Selector4~5_combout )))

	.dataa(\ShiftRight0~22_combout ),
	.datab(\Selector0~9_combout ),
	.datac(\Selector4~5_combout ),
	.datad(\Selector4~3_combout ),
	.cin(gnd),
	.combout(\Selector4~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~6 .lut_mask = 16'hFF40;
defparam \Selector4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N20
cycloneive_lcell_comb \Selector5~2 (
// Equation(s):
// \Selector5~2_combout  = (\portB~13_combout  & ((\Selector0~5_combout ) # ((Mux5 & \Selector0~6_combout ))))

	.dataa(\Selector0~5_combout ),
	.datab(Mux5),
	.datac(\Selector0~6_combout ),
	.datad(portB5),
	.cin(gnd),
	.combout(\Selector5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~2 .lut_mask = 16'hEA00;
defparam \Selector5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N26
cycloneive_lcell_comb \Selector5~3 (
// Equation(s):
// \Selector5~3_combout  = (\Selector5~2_combout ) # ((!Mux5 & (\Selector0~7_combout  & !\portB~13_combout )))

	.dataa(Mux5),
	.datab(\Selector5~2_combout ),
	.datac(\Selector0~7_combout ),
	.datad(portB5),
	.cin(gnd),
	.combout(\Selector5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~3 .lut_mask = 16'hCCDC;
defparam \Selector5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N8
cycloneive_lcell_comb \Selector5~4 (
// Equation(s):
// \Selector5~4_combout  = (\Selector5~3_combout ) # ((\Selector0~11_combout  & (Mux5 $ (\portB~13_combout ))))

	.dataa(\Selector0~11_combout ),
	.datab(Mux5),
	.datac(\Selector5~3_combout ),
	.datad(portB5),
	.cin(gnd),
	.combout(\Selector5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~4 .lut_mask = 16'hF2F8;
defparam \Selector5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N6
cycloneive_lcell_comb \ShiftLeft0~92 (
// Equation(s):
// \ShiftLeft0~92_combout  = (!Mux292 & ((Mux28 & ((\ShiftLeft0~53_combout ))) # (!Mux28 & (\ShiftLeft0~77_combout ))))

	.dataa(Mux292),
	.datab(Mux28),
	.datac(\ShiftLeft0~77_combout ),
	.datad(\ShiftLeft0~53_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~92_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~92 .lut_mask = 16'h5410;
defparam \ShiftLeft0~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N0
cycloneive_lcell_comb \ShiftLeft0~93 (
// Equation(s):
// \ShiftLeft0~93_combout  = (\ShiftLeft0~92_combout ) # ((\Selector7~19_combout  & \ShiftLeft0~73_combout ))

	.dataa(gnd),
	.datab(\Selector7~19_combout ),
	.datac(\ShiftLeft0~73_combout ),
	.datad(\ShiftLeft0~92_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~93_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~93 .lut_mask = 16'hFFC0;
defparam \ShiftLeft0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N18
cycloneive_lcell_comb \ShiftLeft0~86 (
// Equation(s):
// \ShiftLeft0~86_combout  = (\ShiftRight0~122_combout  & ((\portB~25_combout ) # ((\portB~21_combout  & \ShiftRight0~123_combout )))) # (!\ShiftRight0~122_combout  & (((\portB~21_combout  & \ShiftRight0~123_combout ))))

	.dataa(\ShiftRight0~122_combout ),
	.datab(portB11),
	.datac(portB9),
	.datad(\ShiftRight0~123_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~86 .lut_mask = 16'hF888;
defparam \ShiftLeft0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N24
cycloneive_lcell_comb \ShiftLeft0~85 (
// Equation(s):
// \ShiftLeft0~85_combout  = (Mux312 & ((Mux302 & ((\portB~27_combout ))) # (!Mux302 & (\portB~23_combout ))))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB10),
	.datad(portB12),
	.cin(gnd),
	.combout(\ShiftLeft0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~85 .lut_mask = 16'hC840;
defparam \ShiftLeft0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N4
cycloneive_lcell_comb \ShiftLeft0~87 (
// Equation(s):
// \ShiftLeft0~87_combout  = (\ShiftLeft0~86_combout ) # (\ShiftLeft0~85_combout )

	.dataa(gnd),
	.datab(\ShiftLeft0~86_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~85_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~87 .lut_mask = 16'hFFCC;
defparam \ShiftLeft0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N30
cycloneive_lcell_comb \ShiftLeft0~82 (
// Equation(s):
// \ShiftLeft0~82_combout  = (Mux312 & ((Mux302 & ((\portB~35_combout ))) # (!Mux302 & (\portB~31_combout ))))

	.dataa(portB14),
	.datab(portB16),
	.datac(Mux302),
	.datad(Mux312),
	.cin(gnd),
	.combout(\ShiftLeft0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~82 .lut_mask = 16'hCA00;
defparam \ShiftLeft0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N12
cycloneive_lcell_comb \ShiftLeft0~83 (
// Equation(s):
// \ShiftLeft0~83_combout  = (\portB~29_combout  & ((\ShiftRight0~123_combout ) # ((\portB~33_combout  & \ShiftRight0~122_combout )))) # (!\portB~29_combout  & (\portB~33_combout  & (\ShiftRight0~122_combout )))

	.dataa(portB13),
	.datab(portB15),
	.datac(\ShiftRight0~122_combout ),
	.datad(\ShiftRight0~123_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~83 .lut_mask = 16'hEAC0;
defparam \ShiftLeft0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N22
cycloneive_lcell_comb \ShiftLeft0~84 (
// Equation(s):
// \ShiftLeft0~84_combout  = (\ShiftLeft0~82_combout ) # (\ShiftLeft0~83_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftLeft0~82_combout ),
	.datad(\ShiftLeft0~83_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~84 .lut_mask = 16'hFFF0;
defparam \ShiftLeft0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N26
cycloneive_lcell_comb \ShiftLeft0~91 (
// Equation(s):
// \ShiftLeft0~91_combout  = (Mux292 & ((\ShiftLeft0~78_combout ) # ((\ShiftLeft0~79_combout )))) # (!Mux292 & (((\ShiftLeft0~84_combout ))))

	.dataa(Mux292),
	.datab(\ShiftLeft0~78_combout ),
	.datac(\ShiftLeft0~79_combout ),
	.datad(\ShiftLeft0~84_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~91_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~91 .lut_mask = 16'hFDA8;
defparam \ShiftLeft0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N12
cycloneive_lcell_comb \Selector5~5 (
// Equation(s):
// \Selector5~5_combout  = (\Selector7~10_combout  & (\Selector7~18_combout )) # (!\Selector7~10_combout  & ((\Selector7~18_combout  & (\ShiftLeft0~91_combout )) # (!\Selector7~18_combout  & ((\ShiftLeft0~81_combout )))))

	.dataa(\Selector7~10_combout ),
	.datab(\Selector7~18_combout ),
	.datac(\ShiftLeft0~91_combout ),
	.datad(\ShiftLeft0~81_combout ),
	.cin(gnd),
	.combout(\Selector5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~5 .lut_mask = 16'hD9C8;
defparam \Selector5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N2
cycloneive_lcell_comb \Selector5~6 (
// Equation(s):
// \Selector5~6_combout  = (\Selector7~10_combout  & ((\Selector5~5_combout  & (\ShiftLeft0~93_combout )) # (!\Selector5~5_combout  & ((\ShiftLeft0~87_combout ))))) # (!\Selector7~10_combout  & (((\Selector5~5_combout ))))

	.dataa(\Selector7~10_combout ),
	.datab(\ShiftLeft0~93_combout ),
	.datac(\ShiftLeft0~87_combout ),
	.datad(\Selector5~5_combout ),
	.cin(gnd),
	.combout(\Selector5~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~6 .lut_mask = 16'hDDA0;
defparam \Selector5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N24
cycloneive_lcell_comb \Selector5~0 (
// Equation(s):
// \Selector5~0_combout  = (\Selector0~10_combout  & ((\Add0~52_combout ) # ((\Selector0~8_combout  & \Add1~52_combout )))) # (!\Selector0~10_combout  & (\Selector0~8_combout  & (\Add1~52_combout )))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~8_combout ),
	.datac(\Add1~52_combout ),
	.datad(\Add0~52_combout ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~0 .lut_mask = 16'hEAC0;
defparam \Selector5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N2
cycloneive_lcell_comb \Selector5~1 (
// Equation(s):
// \Selector5~1_combout  = (\Selector5~0_combout ) # ((Mux5 & \Selector0~5_combout ))

	.dataa(Mux5),
	.datab(gnd),
	.datac(\Selector0~5_combout ),
	.datad(\Selector5~0_combout ),
	.cin(gnd),
	.combout(\Selector5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~1 .lut_mask = 16'hFFA0;
defparam \Selector5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N12
cycloneive_lcell_comb \ShiftLeft0~23 (
// Equation(s):
// \ShiftLeft0~23_combout  = (\ShiftLeft0~21_combout ) # (\ShiftLeft0~22_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftLeft0~21_combout ),
	.datad(\ShiftLeft0~22_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~23 .lut_mask = 16'hFFF0;
defparam \ShiftLeft0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N20
cycloneive_lcell_comb \Selector12~0 (
// Equation(s):
// \Selector12~0_combout  = (\Selector0~22_combout  & ((Mux292 & (\ShiftLeft0~23_combout )) # (!Mux292 & ((\ShiftLeft0~26_combout )))))

	.dataa(Mux292),
	.datab(\ShiftLeft0~23_combout ),
	.datac(\Selector0~22_combout ),
	.datad(\ShiftLeft0~26_combout ),
	.cin(gnd),
	.combout(\Selector12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~0 .lut_mask = 16'hD080;
defparam \Selector12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N18
cycloneive_lcell_comb \Selector12~1 (
// Equation(s):
// \Selector12~1_combout  = (\Selector12~0_combout ) # ((\Selector1~11_combout  & (\ShiftLeft0~20_combout  & \ShiftRight0~124_combout )))

	.dataa(\Selector1~11_combout ),
	.datab(\ShiftLeft0~20_combout ),
	.datac(\ShiftRight0~124_combout ),
	.datad(\Selector12~0_combout ),
	.cin(gnd),
	.combout(\Selector12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~1 .lut_mask = 16'hFF80;
defparam \Selector12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N4
cycloneive_lcell_comb \ShiftLeft0~10 (
// Equation(s):
// \ShiftLeft0~10_combout  = (\ShiftLeft0~9_combout ) # (\ShiftLeft0~8_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftLeft0~9_combout ),
	.datad(\ShiftLeft0~8_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~10_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~10 .lut_mask = 16'hFFF0;
defparam \ShiftLeft0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N14
cycloneive_lcell_comb \ShiftLeft0~28 (
// Equation(s):
// \ShiftLeft0~28_combout  = (\ShiftRight0~122_combout  & ((\portB~39_combout ) # ((\portB~35_combout  & \ShiftRight0~123_combout )))) # (!\ShiftRight0~122_combout  & (\portB~35_combout  & ((\ShiftRight0~123_combout ))))

	.dataa(\ShiftRight0~122_combout ),
	.datab(portB16),
	.datac(portB18),
	.datad(\ShiftRight0~123_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~28 .lut_mask = 16'hECA0;
defparam \ShiftLeft0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N20
cycloneive_lcell_comb \ShiftLeft0~27 (
// Equation(s):
// \ShiftLeft0~27_combout  = (Mux312 & ((Mux302 & ((\portB~41_combout ))) # (!Mux302 & (\portB~37_combout ))))

	.dataa(portB17),
	.datab(Mux302),
	.datac(Mux312),
	.datad(portB19),
	.cin(gnd),
	.combout(\ShiftLeft0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~27 .lut_mask = 16'hE020;
defparam \ShiftLeft0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N18
cycloneive_lcell_comb \ShiftLeft0~88 (
// Equation(s):
// \ShiftLeft0~88_combout  = (Mux292 & (((\ShiftLeft0~28_combout ) # (\ShiftLeft0~27_combout )))) # (!Mux292 & (\ShiftLeft0~10_combout ))

	.dataa(Mux292),
	.datab(\ShiftLeft0~10_combout ),
	.datac(\ShiftLeft0~28_combout ),
	.datad(\ShiftLeft0~27_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~88 .lut_mask = 16'hEEE4;
defparam \ShiftLeft0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N28
cycloneive_lcell_comb \Selector12~2 (
// Equation(s):
// \Selector12~2_combout  = (\Selector0~14_combout  & ((\Add1~38_combout ) # ((\Selector0~31_combout  & \Add0~38_combout )))) # (!\Selector0~14_combout  & (\Selector0~31_combout  & ((\Add0~38_combout ))))

	.dataa(\Selector0~14_combout ),
	.datab(\Selector0~31_combout ),
	.datac(\Add1~38_combout ),
	.datad(\Add0~38_combout ),
	.cin(gnd),
	.combout(\Selector12~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~2 .lut_mask = 16'hECA0;
defparam \Selector12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N0
cycloneive_lcell_comb \Selector12~6 (
// Equation(s):
// \Selector12~6_combout  = (\Selector12~5_combout ) # ((\Selector12~2_combout ) # ((\Selector0~17_combout  & Mux12)))

	.dataa(\Selector12~5_combout ),
	.datab(\Selector0~17_combout ),
	.datac(Mux12),
	.datad(\Selector12~2_combout ),
	.cin(gnd),
	.combout(\Selector12~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~6 .lut_mask = 16'hFFEA;
defparam \Selector12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N22
cycloneive_lcell_comb \Selector12~7 (
// Equation(s):
// \Selector12~7_combout  = (\Selector12~6_combout ) # ((!cuifALUOP_0 & (\ShiftLeft0~88_combout  & \Selector16~0_combout )))

	.dataa(cuifALUOP_0),
	.datab(\ShiftLeft0~88_combout ),
	.datac(\Selector16~0_combout ),
	.datad(\Selector12~6_combout ),
	.cin(gnd),
	.combout(\Selector12~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~7 .lut_mask = 16'hFF40;
defparam \Selector12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N12
cycloneive_lcell_comb \Selector24~6 (
// Equation(s):
// \Selector24~6_combout  = (\portB~51_combout  & ((\Selector0~5_combout ) # ((\Selector0~6_combout  & Mux242))))

	.dataa(portB24),
	.datab(\Selector0~6_combout ),
	.datac(\Selector0~5_combout ),
	.datad(Mux242),
	.cin(gnd),
	.combout(\Selector24~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~6 .lut_mask = 16'hA8A0;
defparam \Selector24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N30
cycloneive_lcell_comb \Selector24~7 (
// Equation(s):
// \Selector24~7_combout  = (\Selector24~6_combout ) # ((!\portB~51_combout  & (!Mux242 & \Selector0~7_combout )))

	.dataa(portB24),
	.datab(Mux242),
	.datac(\Selector0~7_combout ),
	.datad(\Selector24~6_combout ),
	.cin(gnd),
	.combout(\Selector24~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~7 .lut_mask = 16'hFF10;
defparam \Selector24~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N20
cycloneive_lcell_comb \Selector24~8 (
// Equation(s):
// \Selector24~8_combout  = (\Selector24~7_combout ) # ((\Selector0~11_combout  & (\portB~51_combout  $ (Mux242))))

	.dataa(portB24),
	.datab(\Selector0~11_combout ),
	.datac(\Selector24~7_combout ),
	.datad(Mux242),
	.cin(gnd),
	.combout(\Selector24~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~8 .lut_mask = 16'hF4F8;
defparam \Selector24~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N10
cycloneive_lcell_comb \Selector24~2 (
// Equation(s):
// \Selector24~2_combout  = (\Selector0~10_combout  & ((\Add0~14_combout ) # ((\Selector0~8_combout  & \Add1~14_combout )))) # (!\Selector0~10_combout  & (\Selector0~8_combout  & ((\Add1~14_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~8_combout ),
	.datac(\Add0~14_combout ),
	.datad(\Add1~14_combout ),
	.cin(gnd),
	.combout(\Selector24~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~2 .lut_mask = 16'hECA0;
defparam \Selector24~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N8
cycloneive_lcell_comb \Selector24~1 (
// Equation(s):
// \Selector24~1_combout  = (\Selector0~5_combout  & ((dcifimemload_25 & (Mux24)) # (!dcifimemload_25 & ((Mux241)))))

	.dataa(dcifimemload_25),
	.datab(Mux24),
	.datac(Mux241),
	.datad(\Selector0~5_combout ),
	.cin(gnd),
	.combout(\Selector24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~1 .lut_mask = 16'hD800;
defparam \Selector24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N24
cycloneive_lcell_comb \ShiftRight0~100 (
// Equation(s):
// \ShiftRight0~100_combout  = (Mux292 & (((\ShiftRight0~73_combout ) # (\ShiftRight0~72_combout )))) # (!Mux292 & (\ShiftRight0~61_combout ))

	.dataa(Mux292),
	.datab(\ShiftRight0~61_combout ),
	.datac(\ShiftRight0~73_combout ),
	.datad(\ShiftRight0~72_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~100_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~100 .lut_mask = 16'hEEE4;
defparam \ShiftRight0~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N4
cycloneive_lcell_comb \Selector24~3 (
// Equation(s):
// \Selector24~3_combout  = (\Selector7~18_combout  & (((\Selector7~10_combout )))) # (!\Selector7~18_combout  & ((\Selector7~10_combout  & (\ShiftRight0~101_combout )) # (!\Selector7~10_combout  & ((\ShiftRight0~58_combout )))))

	.dataa(\ShiftRight0~101_combout ),
	.datab(\Selector7~18_combout ),
	.datac(\Selector7~10_combout ),
	.datad(\ShiftRight0~58_combout ),
	.cin(gnd),
	.combout(\Selector24~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~3 .lut_mask = 16'hE3E0;
defparam \Selector24~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N8
cycloneive_lcell_comb \ShiftRight0~65 (
// Equation(s):
// \ShiftRight0~65_combout  = (\ShiftRight0~123_combout  & \portB~3_combout )

	.dataa(gnd),
	.datab(\ShiftRight0~123_combout ),
	.datac(gnd),
	.datad(portB),
	.cin(gnd),
	.combout(\ShiftRight0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~65 .lut_mask = 16'hCC00;
defparam \ShiftRight0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N6
cycloneive_lcell_comb \ShiftRight0~102 (
// Equation(s):
// \ShiftRight0~102_combout  = (Mux292 & (!Mux28 & ((\ShiftRight0~68_combout )))) # (!Mux292 & (Mux28 & (\ShiftRight0~65_combout )))

	.dataa(Mux292),
	.datab(Mux28),
	.datac(\ShiftRight0~65_combout ),
	.datad(\ShiftRight0~68_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~102_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~102 .lut_mask = 16'h6240;
defparam \ShiftRight0~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N24
cycloneive_lcell_comb \ShiftRight0~103 (
// Equation(s):
// \ShiftRight0~103_combout  = (\ShiftRight0~102_combout ) # ((\ShiftRight0~124_combout  & ((\ShiftRight0~70_combout ) # (\ShiftRight0~69_combout ))))

	.dataa(\ShiftRight0~124_combout ),
	.datab(\ShiftRight0~70_combout ),
	.datac(\ShiftRight0~69_combout ),
	.datad(\ShiftRight0~102_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~103_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~103 .lut_mask = 16'hFFA8;
defparam \ShiftRight0~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N24
cycloneive_lcell_comb \Selector24~4 (
// Equation(s):
// \Selector24~4_combout  = (\Selector7~18_combout  & ((\Selector24~3_combout  & ((\ShiftRight0~103_combout ))) # (!\Selector24~3_combout  & (\ShiftRight0~100_combout )))) # (!\Selector7~18_combout  & (((\Selector24~3_combout ))))

	.dataa(\Selector7~18_combout ),
	.datab(\ShiftRight0~100_combout ),
	.datac(\Selector24~3_combout ),
	.datad(\ShiftRight0~103_combout ),
	.cin(gnd),
	.combout(\Selector24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~4 .lut_mask = 16'hF858;
defparam \Selector24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N14
cycloneive_lcell_comb \Selector24~5 (
// Equation(s):
// \Selector24~5_combout  = (\Selector24~2_combout ) # ((\Selector24~1_combout ) # ((Selector24 & \Selector24~4_combout )))

	.dataa(\Selector24~2_combout ),
	.datab(\Selector24~1_combout ),
	.datac(Selector24),
	.datad(\Selector24~4_combout ),
	.cin(gnd),
	.combout(\Selector24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~5 .lut_mask = 16'hFEEE;
defparam \Selector24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N16
cycloneive_lcell_comb \Selector13~0 (
// Equation(s):
// \Selector13~0_combout  = (\Selector0~22_combout  & ((Mux292 & ((\ShiftLeft0~73_combout ))) # (!Mux292 & (\ShiftLeft0~77_combout ))))

	.dataa(\Selector0~22_combout ),
	.datab(\ShiftLeft0~77_combout ),
	.datac(\ShiftLeft0~73_combout ),
	.datad(Mux292),
	.cin(gnd),
	.combout(\Selector13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~0 .lut_mask = 16'hA088;
defparam \Selector13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N14
cycloneive_lcell_comb \Selector13~1 (
// Equation(s):
// \Selector13~1_combout  = (\Selector13~0_combout ) # ((\ShiftRight0~124_combout  & (\Selector1~11_combout  & \ShiftLeft0~53_combout )))

	.dataa(\ShiftRight0~124_combout ),
	.datab(\Selector1~11_combout ),
	.datac(\Selector13~0_combout ),
	.datad(\ShiftLeft0~53_combout ),
	.cin(gnd),
	.combout(\Selector13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~1 .lut_mask = 16'hF8F0;
defparam \Selector13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N12
cycloneive_lcell_comb \Selector13~2 (
// Equation(s):
// \Selector13~2_combout  = (\Selector0~31_combout  & ((\Add0~36_combout ) # ((\Add1~36_combout  & \Selector0~14_combout )))) # (!\Selector0~31_combout  & (\Add1~36_combout  & (\Selector0~14_combout )))

	.dataa(\Selector0~31_combout ),
	.datab(\Add1~36_combout ),
	.datac(\Selector0~14_combout ),
	.datad(\Add0~36_combout ),
	.cin(gnd),
	.combout(\Selector13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~2 .lut_mask = 16'hEAC0;
defparam \Selector13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N0
cycloneive_lcell_comb \Selector13~6 (
// Equation(s):
// \Selector13~6_combout  = (\Selector13~5_combout ) # ((\Selector13~2_combout ) # ((Mux13 & \Selector0~17_combout )))

	.dataa(\Selector13~5_combout ),
	.datab(Mux13),
	.datac(\Selector0~17_combout ),
	.datad(\Selector13~2_combout ),
	.cin(gnd),
	.combout(\Selector13~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~6 .lut_mask = 16'hFFEA;
defparam \Selector13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N22
cycloneive_lcell_comb \Selector13~7 (
// Equation(s):
// \Selector13~7_combout  = (\Selector13~6_combout ) # ((!cuifALUOP_0 & (\Selector16~0_combout  & \ShiftLeft0~91_combout )))

	.dataa(cuifALUOP_0),
	.datab(\Selector16~0_combout ),
	.datac(\ShiftLeft0~91_combout ),
	.datad(\Selector13~6_combout ),
	.cin(gnd),
	.combout(\Selector13~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~7 .lut_mask = 16'hFF40;
defparam \Selector13~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N0
cycloneive_lcell_comb \Selector25~5 (
// Equation(s):
// \Selector25~5_combout  = (\portB~53_combout  & ((\Selector0~5_combout ) # ((Mux252 & \Selector0~6_combout ))))

	.dataa(portB25),
	.datab(Mux252),
	.datac(\Selector0~5_combout ),
	.datad(\Selector0~6_combout ),
	.cin(gnd),
	.combout(\Selector25~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~5 .lut_mask = 16'hA8A0;
defparam \Selector25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N22
cycloneive_lcell_comb \Selector25~6 (
// Equation(s):
// \Selector25~6_combout  = (\Selector25~5_combout ) # ((!\portB~53_combout  & (!Mux252 & \Selector0~7_combout )))

	.dataa(portB25),
	.datab(Mux252),
	.datac(\Selector0~7_combout ),
	.datad(\Selector25~5_combout ),
	.cin(gnd),
	.combout(\Selector25~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~6 .lut_mask = 16'hFF10;
defparam \Selector25~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N8
cycloneive_lcell_comb \Selector25~7 (
// Equation(s):
// \Selector25~7_combout  = (\Selector25~6_combout ) # ((\Selector0~11_combout  & (\portB~53_combout  $ (Mux252))))

	.dataa(portB25),
	.datab(Mux252),
	.datac(\Selector25~6_combout ),
	.datad(\Selector0~11_combout ),
	.cin(gnd),
	.combout(\Selector25~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~7 .lut_mask = 16'hF6F0;
defparam \Selector25~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N26
cycloneive_lcell_comb \Selector25~0 (
// Equation(s):
// \Selector25~0_combout  = (\Selector0~5_combout  & ((dcifimemload_25 & (Mux25)) # (!dcifimemload_25 & ((Mux251)))))

	.dataa(\Selector0~5_combout ),
	.datab(dcifimemload_25),
	.datac(Mux25),
	.datad(Mux251),
	.cin(gnd),
	.combout(\Selector25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~0 .lut_mask = 16'hA280;
defparam \Selector25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N26
cycloneive_lcell_comb \Selector0~10 (
// Equation(s):
// \Selector0~10_combout  = (cuifALUOP_1 & (!cuifALUOP_3 & (!cuifALUOP_0 & !cuifALUOP_2)))

	.dataa(cuifALUOP_1),
	.datab(cuifALUOP_3),
	.datac(cuifALUOP_0),
	.datad(cuifALUOP_2),
	.cin(gnd),
	.combout(\Selector0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~10 .lut_mask = 16'h0002;
defparam \Selector0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N4
cycloneive_lcell_comb \Selector25~1 (
// Equation(s):
// \Selector25~1_combout  = (\Selector0~8_combout  & ((\Add1~12_combout ) # ((\Selector0~10_combout  & \Add0~12_combout )))) # (!\Selector0~8_combout  & (\Selector0~10_combout  & (\Add0~12_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~10_combout ),
	.datac(\Add0~12_combout ),
	.datad(\Add1~12_combout ),
	.cin(gnd),
	.combout(\Selector25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~1 .lut_mask = 16'hEAC0;
defparam \Selector25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N24
cycloneive_lcell_comb \ShiftRight0~105 (
// Equation(s):
// \ShiftRight0~105_combout  = (Mux292 & ((\ShiftRight0~88_combout ) # ((\ShiftRight0~89_combout )))) # (!Mux292 & (((\ShiftRight0~78_combout ))))

	.dataa(\ShiftRight0~88_combout ),
	.datab(\ShiftRight0~89_combout ),
	.datac(Mux292),
	.datad(\ShiftRight0~78_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~105_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~105 .lut_mask = 16'hEFE0;
defparam \ShiftRight0~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N8
cycloneive_lcell_comb \Selector25~2 (
// Equation(s):
// \Selector25~2_combout  = (\Selector7~18_combout  & ((\Selector7~10_combout ) # ((\ShiftRight0~105_combout )))) # (!\Selector7~18_combout  & (!\Selector7~10_combout  & (\ShiftRight0~76_combout )))

	.dataa(\Selector7~18_combout ),
	.datab(\Selector7~10_combout ),
	.datac(\ShiftRight0~76_combout ),
	.datad(\ShiftRight0~105_combout ),
	.cin(gnd),
	.combout(\Selector25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~2 .lut_mask = 16'hBA98;
defparam \Selector25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N14
cycloneive_lcell_comb \ShiftRight0~107 (
// Equation(s):
// \ShiftRight0~107_combout  = (\ShiftRight0~106_combout  & ((Mux28) # ((\Selector7~19_combout  & \ShiftRight0~84_combout )))) # (!\ShiftRight0~106_combout  & (((\Selector7~19_combout  & \ShiftRight0~84_combout ))))

	.dataa(\ShiftRight0~106_combout ),
	.datab(Mux28),
	.datac(\Selector7~19_combout ),
	.datad(\ShiftRight0~84_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~107_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~107 .lut_mask = 16'hF888;
defparam \ShiftRight0~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N10
cycloneive_lcell_comb \ShiftRight0~108 (
// Equation(s):
// \ShiftRight0~108_combout  = (\ShiftRight0~107_combout ) # ((\ShiftRight0~124_combout  & \ShiftRight0~87_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~124_combout ),
	.datac(\ShiftRight0~107_combout ),
	.datad(\ShiftRight0~87_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~108_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~108 .lut_mask = 16'hFCF0;
defparam \ShiftRight0~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N16
cycloneive_lcell_comb \Selector25~3 (
// Equation(s):
// \Selector25~3_combout  = (\Selector7~10_combout  & ((\Selector25~2_combout  & ((\ShiftRight0~108_combout ))) # (!\Selector25~2_combout  & (\ShiftRight0~104_combout )))) # (!\Selector7~10_combout  & (((\Selector25~2_combout ))))

	.dataa(\ShiftRight0~104_combout ),
	.datab(\Selector7~10_combout ),
	.datac(\Selector25~2_combout ),
	.datad(\ShiftRight0~108_combout ),
	.cin(gnd),
	.combout(\Selector25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~3 .lut_mask = 16'hF838;
defparam \Selector25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N2
cycloneive_lcell_comb \Selector25~4 (
// Equation(s):
// \Selector25~4_combout  = (\Selector25~0_combout ) # ((\Selector25~1_combout ) # ((Selector24 & \Selector25~3_combout )))

	.dataa(Selector24),
	.datab(\Selector25~0_combout ),
	.datac(\Selector25~1_combout ),
	.datad(\Selector25~3_combout ),
	.cin(gnd),
	.combout(\Selector25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~4 .lut_mask = 16'hFEFC;
defparam \Selector25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N12
cycloneive_lcell_comb \Selector1~25 (
// Equation(s):
// \Selector1~25_combout  = (Mux302) # ((dcifimemload_25 & ((Mux29))) # (!dcifimemload_25 & (Mux291)))

	.dataa(dcifimemload_25),
	.datab(Mux291),
	.datac(Mux302),
	.datad(Mux29),
	.cin(gnd),
	.combout(\Selector1~25_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~25 .lut_mask = 16'hFEF4;
defparam \Selector1~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N30
cycloneive_lcell_comb \ShiftLeft0~94 (
// Equation(s):
// \ShiftLeft0~94_combout  = (!\Selector1~25_combout  & ((Mux312 & (\portB~65_combout )) # (!Mux312 & ((\portB~63_combout )))))

	.dataa(portB31),
	.datab(\Selector1~25_combout ),
	.datac(portB30),
	.datad(Mux312),
	.cin(gnd),
	.combout(\ShiftLeft0~94_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~94 .lut_mask = 16'h2230;
defparam \ShiftLeft0~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N4
cycloneive_lcell_comb \Selector14~0 (
// Equation(s):
// \Selector14~0_combout  = (Mux292 & ((\ShiftLeft0~55_combout ) # ((\ShiftLeft0~54_combout )))) # (!Mux292 & (((\ShiftLeft0~59_combout ))))

	.dataa(\ShiftLeft0~55_combout ),
	.datab(Mux292),
	.datac(\ShiftLeft0~54_combout ),
	.datad(\ShiftLeft0~59_combout ),
	.cin(gnd),
	.combout(\Selector14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~0 .lut_mask = 16'hFBC8;
defparam \Selector14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N24
cycloneive_lcell_comb \Selector14~3 (
// Equation(s):
// \Selector14~3_combout  = (\portB~31_combout  & ((\Selector0~17_combout ) # ((\Selector0~18_combout  & Mux14))))

	.dataa(\Selector0~17_combout ),
	.datab(portB14),
	.datac(\Selector0~18_combout ),
	.datad(Mux14),
	.cin(gnd),
	.combout(\Selector14~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~3 .lut_mask = 16'hC888;
defparam \Selector14~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N26
cycloneive_lcell_comb \Selector14~4 (
// Equation(s):
// \Selector14~4_combout  = (\Selector14~3_combout ) # ((\Selector0~27_combout  & (!Mux14 & !\portB~31_combout )))

	.dataa(\Selector0~27_combout ),
	.datab(\Selector14~3_combout ),
	.datac(Mux14),
	.datad(portB14),
	.cin(gnd),
	.combout(\Selector14~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~4 .lut_mask = 16'hCCCE;
defparam \Selector14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N4
cycloneive_lcell_comb \Selector14~5 (
// Equation(s):
// \Selector14~5_combout  = (\Selector14~4_combout ) # ((\Selector0~15_combout  & (\portB~31_combout  $ (Mux14))))

	.dataa(\Selector14~4_combout ),
	.datab(portB14),
	.datac(\Selector0~15_combout ),
	.datad(Mux14),
	.cin(gnd),
	.combout(\Selector14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~5 .lut_mask = 16'hBAEA;
defparam \Selector14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N6
cycloneive_lcell_comb \Selector14~2 (
// Equation(s):
// \Selector14~2_combout  = (\Selector0~31_combout  & ((\Add0~34_combout ) # ((\Selector0~14_combout  & \Add1~34_combout )))) # (!\Selector0~31_combout  & (\Selector0~14_combout  & (\Add1~34_combout )))

	.dataa(\Selector0~31_combout ),
	.datab(\Selector0~14_combout ),
	.datac(\Add1~34_combout ),
	.datad(\Add0~34_combout ),
	.cin(gnd),
	.combout(\Selector14~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~2 .lut_mask = 16'hEAC0;
defparam \Selector14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N22
cycloneive_lcell_comb \ShiftLeft0~64 (
// Equation(s):
// \ShiftLeft0~64_combout  = (\ShiftLeft0~63_combout ) # (\ShiftLeft0~62_combout )

	.dataa(\ShiftLeft0~63_combout ),
	.datab(gnd),
	.datac(\ShiftLeft0~62_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~64 .lut_mask = 16'hFAFA;
defparam \ShiftLeft0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N8
cycloneive_lcell_comb \ShiftLeft0~95 (
// Equation(s):
// \ShiftLeft0~95_combout  = (Mux292 & ((\ShiftLeft0~61_combout ) # ((\ShiftLeft0~60_combout )))) # (!Mux292 & (((\ShiftLeft0~64_combout ))))

	.dataa(\ShiftLeft0~61_combout ),
	.datab(Mux292),
	.datac(\ShiftLeft0~64_combout ),
	.datad(\ShiftLeft0~60_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~95_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~95 .lut_mask = 16'hFCB8;
defparam \ShiftLeft0~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N2
cycloneive_lcell_comb \ShiftRight0~92 (
// Equation(s):
// \ShiftRight0~92_combout  = (Mux302 & ((Mux312 & (\portB~9_combout )) # (!Mux312 & ((\portB~11_combout )))))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB3),
	.datad(portB4),
	.cin(gnd),
	.combout(\ShiftRight0~92_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~92 .lut_mask = 16'hA280;
defparam \ShiftRight0~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N20
cycloneive_lcell_comb \ShiftRight0~91 (
// Equation(s):
// \ShiftRight0~91_combout  = (!Mux302 & (Mux312 & \portB~13_combout ))

	.dataa(Mux302),
	.datab(gnd),
	.datac(Mux312),
	.datad(portB5),
	.cin(gnd),
	.combout(\ShiftRight0~91_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~91 .lut_mask = 16'h5000;
defparam \ShiftRight0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N12
cycloneive_lcell_comb \ShiftRight0~93 (
// Equation(s):
// \ShiftRight0~93_combout  = (\ShiftRight0~92_combout ) # ((\ShiftRight0~91_combout ) # ((\ShiftRight0~123_combout  & \portB~15_combout )))

	.dataa(\ShiftRight0~123_combout ),
	.datab(\ShiftRight0~92_combout ),
	.datac(portB6),
	.datad(\ShiftRight0~91_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~93_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~93 .lut_mask = 16'hFFEC;
defparam \ShiftRight0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N2
cycloneive_lcell_comb \ShiftRight0~109 (
// Equation(s):
// \ShiftRight0~109_combout  = (Mux292 & (\ShiftRight0~98_combout )) # (!Mux292 & ((\ShiftRight0~93_combout )))

	.dataa(\ShiftRight0~98_combout ),
	.datab(gnd),
	.datac(\ShiftRight0~93_combout ),
	.datad(Mux292),
	.cin(gnd),
	.combout(\ShiftRight0~109_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~109 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N8
cycloneive_lcell_comb \ShiftRight0~110 (
// Equation(s):
// \ShiftRight0~110_combout  = (Mux312 & ((\portB~25_combout ) # ((!Mux302)))) # (!Mux312 & (((\portB~27_combout  & Mux302))))

	.dataa(Mux312),
	.datab(portB11),
	.datac(portB12),
	.datad(Mux302),
	.cin(gnd),
	.combout(\ShiftRight0~110_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~110 .lut_mask = 16'hD8AA;
defparam \ShiftRight0~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N30
cycloneive_lcell_comb \ShiftRight0~111 (
// Equation(s):
// \ShiftRight0~111_combout  = (\ShiftRight0~110_combout  & ((\portB~29_combout ) # ((Mux302)))) # (!\ShiftRight0~110_combout  & (((\portB~31_combout  & !Mux302))))

	.dataa(portB13),
	.datab(\ShiftRight0~110_combout ),
	.datac(portB14),
	.datad(Mux302),
	.cin(gnd),
	.combout(\ShiftRight0~111_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~111 .lut_mask = 16'hCCB8;
defparam \ShiftRight0~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N18
cycloneive_lcell_comb \Selector22~1 (
// Equation(s):
// \Selector22~1_combout  = (Mux292 & ((\ShiftRight0~95_combout ))) # (!Mux292 & (\ShiftRight0~111_combout ))

	.dataa(gnd),
	.datab(Mux292),
	.datac(\ShiftRight0~111_combout ),
	.datad(\ShiftRight0~95_combout ),
	.cin(gnd),
	.combout(\Selector22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~1 .lut_mask = 16'hFC30;
defparam \Selector22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N28
cycloneive_lcell_comb \ShiftRight0~112 (
// Equation(s):
// \ShiftRight0~112_combout  = (Mux28 & (\ShiftRight0~109_combout )) # (!Mux28 & ((\Selector22~1_combout )))

	.dataa(gnd),
	.datab(Mux28),
	.datac(\ShiftRight0~109_combout ),
	.datad(\Selector22~1_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~112_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~112 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~112 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N2
cycloneive_lcell_comb \Selector27~5 (
// Equation(s):
// \Selector27~5_combout  = (\portB~57_combout  & ((\Selector0~5_combout ) # ((Mux272 & \Selector0~6_combout ))))

	.dataa(Mux272),
	.datab(portB27),
	.datac(\Selector0~5_combout ),
	.datad(\Selector0~6_combout ),
	.cin(gnd),
	.combout(\Selector27~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~5 .lut_mask = 16'hC8C0;
defparam \Selector27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N4
cycloneive_lcell_comb \Selector27~6 (
// Equation(s):
// \Selector27~6_combout  = (\Selector27~5_combout ) # ((!\portB~57_combout  & (\Selector0~7_combout  & !Mux272)))

	.dataa(portB27),
	.datab(\Selector0~7_combout ),
	.datac(Mux272),
	.datad(\Selector27~5_combout ),
	.cin(gnd),
	.combout(\Selector27~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~6 .lut_mask = 16'hFF04;
defparam \Selector27~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N22
cycloneive_lcell_comb \Selector27~7 (
// Equation(s):
// \Selector27~7_combout  = (\Selector27~6_combout ) # ((\Selector0~11_combout  & (Mux272 $ (\portB~57_combout ))))

	.dataa(Mux272),
	.datab(portB27),
	.datac(\Selector27~6_combout ),
	.datad(\Selector0~11_combout ),
	.cin(gnd),
	.combout(\Selector27~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~7 .lut_mask = 16'hF6F0;
defparam \Selector27~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N28
cycloneive_lcell_comb \Selector27~0 (
// Equation(s):
// \Selector27~0_combout  = (\Selector0~10_combout  & ((\Add0~8_combout ) # ((\Selector0~8_combout  & \Add1~8_combout )))) # (!\Selector0~10_combout  & (\Selector0~8_combout  & ((\Add1~8_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~8_combout ),
	.datac(\Add0~8_combout ),
	.datad(\Add1~8_combout ),
	.cin(gnd),
	.combout(\Selector27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~0 .lut_mask = 16'hECA0;
defparam \Selector27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N2
cycloneive_lcell_comb \Selector27~1 (
// Equation(s):
// \Selector27~1_combout  = (\Selector27~0_combout ) # ((\Selector0~5_combout  & Mux272))

	.dataa(\Selector0~5_combout ),
	.datab(gnd),
	.datac(Mux272),
	.datad(\Selector27~0_combout ),
	.cin(gnd),
	.combout(\Selector27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~1 .lut_mask = 16'hFFA0;
defparam \Selector27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N12
cycloneive_lcell_comb \Selector27~3 (
// Equation(s):
// \Selector27~3_combout  = (\Selector27~2_combout  & (((ShiftRight01)) # (!\Selector7~10_combout ))) # (!\Selector27~2_combout  & (\Selector7~10_combout  & ((\ShiftRight0~48_combout ))))

	.dataa(\Selector27~2_combout ),
	.datab(\Selector7~10_combout ),
	.datac(ShiftRight01),
	.datad(\ShiftRight0~48_combout ),
	.cin(gnd),
	.combout(\Selector27~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~3 .lut_mask = 16'hE6A2;
defparam \Selector27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N22
cycloneive_lcell_comb \Selector27~4 (
// Equation(s):
// \Selector27~4_combout  = (\Selector27~1_combout ) # ((\Selector0~13_combout  & (!\ShiftRight0~22_combout  & \Selector27~3_combout )))

	.dataa(\Selector0~13_combout ),
	.datab(\ShiftRight0~22_combout ),
	.datac(\Selector27~1_combout ),
	.datad(\Selector27~3_combout ),
	.cin(gnd),
	.combout(\Selector27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~4 .lut_mask = 16'hF2F0;
defparam \Selector27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N10
cycloneive_lcell_comb \Selector8~1 (
// Equation(s):
// \Selector8~1_combout  = (Mux292 & (\ShiftLeft0~26_combout )) # (!Mux292 & (((\ShiftLeft0~28_combout ) # (\ShiftLeft0~27_combout ))))

	.dataa(Mux292),
	.datab(\ShiftLeft0~26_combout ),
	.datac(\ShiftLeft0~28_combout ),
	.datad(\ShiftLeft0~27_combout ),
	.cin(gnd),
	.combout(\Selector8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~1 .lut_mask = 16'hDDD8;
defparam \Selector8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N26
cycloneive_lcell_comb \ShiftLeft0~96 (
// Equation(s):
// \ShiftLeft0~96_combout  = (Mux28 & ((\ShiftLeft0~101_combout ))) # (!Mux28 & (\Selector8~1_combout ))

	.dataa(\Selector8~1_combout ),
	.datab(\ShiftLeft0~101_combout ),
	.datac(Mux28),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~96_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~96 .lut_mask = 16'hCACA;
defparam \ShiftLeft0~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N12
cycloneive_lcell_comb \Selector16~3 (
// Equation(s):
// \Selector16~3_combout  = (\portB~35_combout  & ((\Selector0~17_combout ) # ((Mux16 & \Selector0~18_combout ))))

	.dataa(portB16),
	.datab(\Selector0~17_combout ),
	.datac(Mux16),
	.datad(\Selector0~18_combout ),
	.cin(gnd),
	.combout(\Selector16~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~3 .lut_mask = 16'hA888;
defparam \Selector16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N2
cycloneive_lcell_comb \Selector16~4 (
// Equation(s):
// \Selector16~4_combout  = (\Selector16~3_combout ) # ((!\portB~35_combout  & (\Selector0~27_combout  & !Mux16)))

	.dataa(portB16),
	.datab(\Selector0~27_combout ),
	.datac(Mux16),
	.datad(\Selector16~3_combout ),
	.cin(gnd),
	.combout(\Selector16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~4 .lut_mask = 16'hFF04;
defparam \Selector16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N4
cycloneive_lcell_comb \Selector16~5 (
// Equation(s):
// \Selector16~5_combout  = (\Selector16~4_combout ) # ((\Selector0~15_combout  & (Mux16 $ (\portB~35_combout ))))

	.dataa(\Selector0~15_combout ),
	.datab(Mux16),
	.datac(portB16),
	.datad(\Selector16~4_combout ),
	.cin(gnd),
	.combout(\Selector16~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~5 .lut_mask = 16'hFF28;
defparam \Selector16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N18
cycloneive_lcell_comb \Selector16~2 (
// Equation(s):
// \Selector16~2_combout  = (\Selector0~14_combout  & ((\Add1~30_combout ) # ((\Selector0~31_combout  & \Add0~30_combout )))) # (!\Selector0~14_combout  & (\Selector0~31_combout  & ((\Add0~30_combout ))))

	.dataa(\Selector0~14_combout ),
	.datab(\Selector0~31_combout ),
	.datac(\Add1~30_combout ),
	.datad(\Add0~30_combout ),
	.cin(gnd),
	.combout(\Selector16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~2 .lut_mask = 16'hECA0;
defparam \Selector16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N30
cycloneive_lcell_comb \Selector16~6 (
// Equation(s):
// \Selector16~6_combout  = (\Selector16~5_combout ) # ((\Selector16~2_combout ) # ((\Selector0~17_combout  & Mux16)))

	.dataa(\Selector0~17_combout ),
	.datab(Mux16),
	.datac(\Selector16~5_combout ),
	.datad(\Selector16~2_combout ),
	.cin(gnd),
	.combout(\Selector16~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~6 .lut_mask = 16'hFFF8;
defparam \Selector16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N26
cycloneive_lcell_comb \Selector16~9 (
// Equation(s):
// \Selector16~9_combout  = (cuifALUOP_0 & \Selector16~0_combout )

	.dataa(cuifALUOP_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\Selector16~0_combout ),
	.cin(gnd),
	.combout(\Selector16~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~9 .lut_mask = 16'hAA00;
defparam \Selector16~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N10
cycloneive_lcell_comb \Selector16~8 (
// Equation(s):
// \Selector16~8_combout  = (!\ShiftRight0~23_combout  & (\portB~3_combout  & Selector22))

	.dataa(\ShiftRight0~23_combout ),
	.datab(portB),
	.datac(gnd),
	.datad(Selector22),
	.cin(gnd),
	.combout(\Selector16~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~8 .lut_mask = 16'h4400;
defparam \Selector16~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N16
cycloneive_lcell_comb \Selector0~35 (
// Equation(s):
// \Selector0~35_combout  = (cuifALUOP_0 & (Mux28 & (\Selector1~8_combout  & !Mux272)))

	.dataa(cuifALUOP_0),
	.datab(Mux28),
	.datac(\Selector1~8_combout ),
	.datad(Mux272),
	.cin(gnd),
	.combout(\Selector0~35_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~35 .lut_mask = 16'h0080;
defparam \Selector0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N28
cycloneive_lcell_comb \Selector16~7 (
// Equation(s):
// \Selector16~7_combout  = (\Selector0~35_combout  & ((Mux292 & (\ShiftRight0~68_combout )) # (!Mux292 & ((\ShiftRight0~71_combout )))))

	.dataa(\ShiftRight0~68_combout ),
	.datab(Mux292),
	.datac(\Selector0~35_combout ),
	.datad(\ShiftRight0~71_combout ),
	.cin(gnd),
	.combout(\Selector16~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~7 .lut_mask = 16'hB080;
defparam \Selector16~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N10
cycloneive_lcell_comb \Selector16~10 (
// Equation(s):
// \Selector16~10_combout  = (\Selector16~8_combout ) # ((\Selector16~7_combout ) # ((\Selector16~9_combout  & \ShiftRight0~100_combout )))

	.dataa(\Selector16~9_combout ),
	.datab(\ShiftRight0~100_combout ),
	.datac(\Selector16~8_combout ),
	.datad(\Selector16~7_combout ),
	.cin(gnd),
	.combout(\Selector16~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~10 .lut_mask = 16'hFFF8;
defparam \Selector16~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N2
cycloneive_lcell_comb \Selector18~0 (
// Equation(s):
// \Selector18~0_combout  = (\Selector0~35_combout  & ((Mux292 & ((\ShiftRight0~93_combout ))) # (!Mux292 & (\ShiftRight0~95_combout ))))

	.dataa(\ShiftRight0~95_combout ),
	.datab(Mux292),
	.datac(\Selector0~35_combout ),
	.datad(\ShiftRight0~93_combout ),
	.cin(gnd),
	.combout(\Selector18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~0 .lut_mask = 16'hE020;
defparam \Selector18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N0
cycloneive_lcell_comb \Selector18~1 (
// Equation(s):
// \Selector18~1_combout  = (\Selector18~0_combout ) # ((\ShiftRight0~98_combout  & (Selector22 & \ShiftRight0~124_combout )))

	.dataa(\ShiftRight0~98_combout ),
	.datab(Selector22),
	.datac(\ShiftRight0~124_combout ),
	.datad(\Selector18~0_combout ),
	.cin(gnd),
	.combout(\Selector18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~1 .lut_mask = 16'hFF80;
defparam \Selector18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N6
cycloneive_lcell_comb \Selector18~2 (
// Equation(s):
// \Selector18~2_combout  = (\Add1~26_combout  & ((\Selector0~14_combout ) # ((\Selector0~31_combout  & \Add0~26_combout )))) # (!\Add1~26_combout  & (\Selector0~31_combout  & ((\Add0~26_combout ))))

	.dataa(\Add1~26_combout ),
	.datab(\Selector0~31_combout ),
	.datac(\Selector0~14_combout ),
	.datad(\Add0~26_combout ),
	.cin(gnd),
	.combout(\Selector18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~2 .lut_mask = 16'hECA0;
defparam \Selector18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N30
cycloneive_lcell_comb \Selector18~6 (
// Equation(s):
// \Selector18~6_combout  = (\Selector18~5_combout ) # ((\Selector18~2_combout ) # ((\Selector0~17_combout  & Mux18)))

	.dataa(\Selector18~5_combout ),
	.datab(\Selector0~17_combout ),
	.datac(Mux18),
	.datad(\Selector18~2_combout ),
	.cin(gnd),
	.combout(\Selector18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~6 .lut_mask = 16'hFFEA;
defparam \Selector18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N0
cycloneive_lcell_comb \ShiftRight0~115 (
// Equation(s):
// \ShiftRight0~115_combout  = (Mux302 & ((Mux312 & ((\portB~33_combout ))) # (!Mux312 & (\portB~35_combout ))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB16),
	.datad(portB15),
	.cin(gnd),
	.combout(\ShiftRight0~115_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~115 .lut_mask = 16'hC840;
defparam \ShiftRight0~115 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N30
cycloneive_lcell_comb \ShiftRight0~114 (
// Equation(s):
// \ShiftRight0~114_combout  = (!Mux302 & ((Mux312 & (\portB~37_combout )) # (!Mux312 & ((\portB~39_combout )))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB17),
	.datad(portB18),
	.cin(gnd),
	.combout(\ShiftRight0~114_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~114 .lut_mask = 16'h3120;
defparam \ShiftRight0~114 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N14
cycloneive_lcell_comb \ShiftRight0~116 (
// Equation(s):
// \ShiftRight0~116_combout  = (Mux292 & (((\ShiftRight0~111_combout )))) # (!Mux292 & ((\ShiftRight0~115_combout ) # ((\ShiftRight0~114_combout ))))

	.dataa(Mux292),
	.datab(\ShiftRight0~115_combout ),
	.datac(\ShiftRight0~114_combout ),
	.datad(\ShiftRight0~111_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~116_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~116 .lut_mask = 16'hFE54;
defparam \ShiftRight0~116 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N4
cycloneive_lcell_comb \Selector18~7 (
// Equation(s):
// \Selector18~7_combout  = (\Selector18~6_combout ) # ((cuifALUOP_0 & (\Selector16~0_combout  & \ShiftRight0~116_combout )))

	.dataa(cuifALUOP_0),
	.datab(\Selector16~0_combout ),
	.datac(\Selector18~6_combout ),
	.datad(\ShiftRight0~116_combout ),
	.cin(gnd),
	.combout(\Selector18~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~7 .lut_mask = 16'hF8F0;
defparam \Selector18~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N8
cycloneive_lcell_comb \ShiftLeft0~97 (
// Equation(s):
// \ShiftLeft0~97_combout  = (Mux28 & (ShiftLeft0)) # (!Mux28 & ((\Selector10~0_combout )))

	.dataa(Mux28),
	.datab(gnd),
	.datac(ShiftLeft0),
	.datad(\Selector10~0_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~97_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~97 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N22
cycloneive_lcell_comb \ShiftLeft0~98 (
// Equation(s):
// \ShiftLeft0~98_combout  = (Mux28 & (\ShiftLeft0~74_combout )) # (!Mux28 & ((\Selector9~0_combout )))

	.dataa(gnd),
	.datab(Mux28),
	.datac(\ShiftLeft0~74_combout ),
	.datad(\Selector9~0_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~98_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~98 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N6
cycloneive_lcell_comb \Selector17~0 (
// Equation(s):
// \Selector17~0_combout  = (Mux292 & (\ShiftRight0~84_combout )) # (!Mux292 & ((\ShiftRight0~87_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~84_combout ),
	.datac(Mux292),
	.datad(\ShiftRight0~87_combout ),
	.cin(gnd),
	.combout(\Selector17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~0 .lut_mask = 16'hCFC0;
defparam \Selector17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N8
cycloneive_lcell_comb \Selector17~1 (
// Equation(s):
// \Selector17~1_combout  = (\Selector0~35_combout  & ((\Selector17~0_combout ) # ((\ShiftRight0~105_combout  & \Selector16~9_combout )))) # (!\Selector0~35_combout  & (\ShiftRight0~105_combout  & ((\Selector16~9_combout ))))

	.dataa(\Selector0~35_combout ),
	.datab(\ShiftRight0~105_combout ),
	.datac(\Selector17~0_combout ),
	.datad(\Selector16~9_combout ),
	.cin(gnd),
	.combout(\Selector17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~1 .lut_mask = 16'hECA0;
defparam \Selector17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N12
cycloneive_lcell_comb \ShiftRight0~106 (
// Equation(s):
// \ShiftRight0~106_combout  = (!\Selector1~25_combout  & ((Mux312 & (\portB~3_combout )) # (!Mux312 & ((\portB~5_combout )))))

	.dataa(Mux312),
	.datab(\Selector1~25_combout ),
	.datac(portB),
	.datad(portB1),
	.cin(gnd),
	.combout(\ShiftRight0~106_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~106 .lut_mask = 16'h3120;
defparam \ShiftRight0~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N18
cycloneive_lcell_comb \Selector17~2 (
// Equation(s):
// \Selector17~2_combout  = (\Selector0~31_combout  & ((\Add0~28_combout ) # ((\Selector0~14_combout  & \Add1~28_combout )))) # (!\Selector0~31_combout  & (\Selector0~14_combout  & (\Add1~28_combout )))

	.dataa(\Selector0~31_combout ),
	.datab(\Selector0~14_combout ),
	.datac(\Add1~28_combout ),
	.datad(\Add0~28_combout ),
	.cin(gnd),
	.combout(\Selector17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~2 .lut_mask = 16'hEAC0;
defparam \Selector17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N14
cycloneive_lcell_comb \Selector17~6 (
// Equation(s):
// \Selector17~6_combout  = (\Selector17~5_combout ) # ((\Selector17~2_combout ) # ((\Selector0~17_combout  & Mux17)))

	.dataa(\Selector17~5_combout ),
	.datab(\Selector0~17_combout ),
	.datac(Mux17),
	.datad(\Selector17~2_combout ),
	.cin(gnd),
	.combout(\Selector17~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~6 .lut_mask = 16'hFFEA;
defparam \Selector17~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N12
cycloneive_lcell_comb \Selector17~7 (
// Equation(s):
// \Selector17~7_combout  = (\Selector17~6_combout ) # ((\ShiftRight0~106_combout  & (!Mux28 & Selector22)))

	.dataa(\ShiftRight0~106_combout ),
	.datab(Mux28),
	.datac(\Selector17~6_combout ),
	.datad(Selector22),
	.cin(gnd),
	.combout(\Selector17~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~7 .lut_mask = 16'hF2F0;
defparam \Selector17~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N26
cycloneive_lcell_comb \Selector6~2 (
// Equation(s):
// \Selector6~2_combout  = (\portB~15_combout  & ((\Selector0~5_combout ) # ((Mux6 & \Selector0~6_combout ))))

	.dataa(Mux6),
	.datab(portB6),
	.datac(\Selector0~5_combout ),
	.datad(\Selector0~6_combout ),
	.cin(gnd),
	.combout(\Selector6~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~2 .lut_mask = 16'hC8C0;
defparam \Selector6~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N22
cycloneive_lcell_comb \Selector6~5 (
// Equation(s):
// \Selector6~5_combout  = (Mux6 & (\Selector0~11_combout  & ((!\portB~15_combout )))) # (!Mux6 & ((\portB~15_combout  & (\Selector0~11_combout )) # (!\portB~15_combout  & ((\Selector0~7_combout )))))

	.dataa(Mux6),
	.datab(\Selector0~11_combout ),
	.datac(\Selector0~7_combout ),
	.datad(portB6),
	.cin(gnd),
	.combout(\Selector6~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~5 .lut_mask = 16'h44D8;
defparam \Selector6~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N6
cycloneive_lcell_comb \Selector6~3 (
// Equation(s):
// \Selector6~3_combout  = (\Selector0~8_combout  & ((\Add1~50_combout ) # ((\Selector0~10_combout  & \Add0~50_combout )))) # (!\Selector0~8_combout  & (\Selector0~10_combout  & ((\Add0~50_combout ))))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~10_combout ),
	.datac(\Add1~50_combout ),
	.datad(\Add0~50_combout ),
	.cin(gnd),
	.combout(\Selector6~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~3 .lut_mask = 16'hECA0;
defparam \Selector6~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N28
cycloneive_lcell_comb \Selector6~4 (
// Equation(s):
// \Selector6~4_combout  = (\Selector6~3_combout ) # ((Mux6 & \Selector0~5_combout ))

	.dataa(Mux6),
	.datab(gnd),
	.datac(\Selector0~5_combout ),
	.datad(\Selector6~3_combout ),
	.cin(gnd),
	.combout(\Selector6~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~4 .lut_mask = 16'hFFA0;
defparam \Selector6~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N30
cycloneive_lcell_comb \Selector6~6 (
// Equation(s):
// \Selector6~6_combout  = (\Selector6~5_combout ) # ((\Selector6~4_combout ) # ((Selector4 & \ShiftRight0~109_combout )))

	.dataa(Selector4),
	.datab(\Selector6~5_combout ),
	.datac(\ShiftRight0~109_combout ),
	.datad(\Selector6~4_combout ),
	.cin(gnd),
	.combout(\Selector6~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~6 .lut_mask = 16'hFFEC;
defparam \Selector6~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N0
cycloneive_lcell_comb \Selector6~0 (
// Equation(s):
// \Selector6~0_combout  = (\Selector7~18_combout  & (\Selector7~10_combout )) # (!\Selector7~18_combout  & ((\Selector7~10_combout  & (\ShiftLeft0~67_combout )) # (!\Selector7~10_combout  & ((\ShiftLeft0~70_combout )))))

	.dataa(\Selector7~18_combout ),
	.datab(\Selector7~10_combout ),
	.datac(\ShiftLeft0~67_combout ),
	.datad(\ShiftLeft0~70_combout ),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~0 .lut_mask = 16'hD9C8;
defparam \Selector6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N12
cycloneive_lcell_comb \ShiftLeft0~99 (
// Equation(s):
// \ShiftLeft0~99_combout  = (Mux28 & ((\ShiftLeft0~94_combout ) # ((\ShiftRight0~124_combout  & \ShiftLeft0~59_combout )))) # (!Mux28 & (\ShiftRight0~124_combout  & ((\ShiftLeft0~59_combout ))))

	.dataa(Mux28),
	.datab(\ShiftRight0~124_combout ),
	.datac(\ShiftLeft0~94_combout ),
	.datad(\ShiftLeft0~59_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~99_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~99 .lut_mask = 16'hECA0;
defparam \ShiftLeft0~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N18
cycloneive_lcell_comb \ShiftLeft0~100 (
// Equation(s):
// \ShiftLeft0~100_combout  = (\ShiftLeft0~99_combout ) # ((\Selector7~19_combout  & ((\ShiftLeft0~55_combout ) # (\ShiftLeft0~54_combout ))))

	.dataa(\ShiftLeft0~55_combout ),
	.datab(\Selector7~19_combout ),
	.datac(\ShiftLeft0~54_combout ),
	.datad(\ShiftLeft0~99_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~100_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~100 .lut_mask = 16'hFFC8;
defparam \ShiftLeft0~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N12
cycloneive_lcell_comb \Selector6~1 (
// Equation(s):
// \Selector6~1_combout  = (\Selector7~18_combout  & ((\Selector6~0_combout  & ((\ShiftLeft0~100_combout ))) # (!\Selector6~0_combout  & (\ShiftLeft0~95_combout )))) # (!\Selector7~18_combout  & (\Selector6~0_combout ))

	.dataa(\Selector7~18_combout ),
	.datab(\Selector6~0_combout ),
	.datac(\ShiftLeft0~95_combout ),
	.datad(\ShiftLeft0~100_combout ),
	.cin(gnd),
	.combout(\Selector6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~1 .lut_mask = 16'hEC64;
defparam \Selector6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N18
cycloneive_lcell_comb \Selector26~0 (
// Equation(s):
// \Selector26~0_combout  = (\Selector0~10_combout  & ((\Add0~10_combout ) # ((\Selector0~8_combout  & \Add1~10_combout )))) # (!\Selector0~10_combout  & (((\Selector0~8_combout  & \Add1~10_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(\Add0~10_combout ),
	.datac(\Selector0~8_combout ),
	.datad(\Add1~10_combout ),
	.cin(gnd),
	.combout(\Selector26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~0 .lut_mask = 16'hF888;
defparam \Selector26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N4
cycloneive_lcell_comb \Selector26~1 (
// Equation(s):
// \Selector26~1_combout  = (\Selector26~0_combout ) # ((\Selector0~5_combout  & Mux26))

	.dataa(\Selector0~5_combout ),
	.datab(gnd),
	.datac(Mux26),
	.datad(\Selector26~0_combout ),
	.cin(gnd),
	.combout(\Selector26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~1 .lut_mask = 16'hFFA0;
defparam \Selector26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N30
cycloneive_lcell_comb \Selector26~2 (
// Equation(s):
// \Selector26~2_combout  = (\portB~55_combout  & ((\Selector0~5_combout ) # ((\Selector0~6_combout  & Mux26))))

	.dataa(portB26),
	.datab(\Selector0~6_combout ),
	.datac(Mux26),
	.datad(\Selector0~5_combout ),
	.cin(gnd),
	.combout(\Selector26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~2 .lut_mask = 16'hAA80;
defparam \Selector26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N8
cycloneive_lcell_comb \Selector26~3 (
// Equation(s):
// \Selector26~3_combout  = (\Selector26~2_combout ) # ((\Selector0~7_combout  & (!Mux26 & !\portB~55_combout )))

	.dataa(\Selector0~7_combout ),
	.datab(Mux26),
	.datac(\Selector26~2_combout ),
	.datad(portB26),
	.cin(gnd),
	.combout(\Selector26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~3 .lut_mask = 16'hF0F2;
defparam \Selector26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N22
cycloneive_lcell_comb \Selector26~4 (
// Equation(s):
// \Selector26~4_combout  = (\Selector26~3_combout ) # ((\Selector0~11_combout  & (Mux26 $ (\portB~55_combout ))))

	.dataa(Mux26),
	.datab(\Selector26~3_combout ),
	.datac(\Selector0~11_combout ),
	.datad(portB26),
	.cin(gnd),
	.combout(\Selector26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~4 .lut_mask = 16'hDCEC;
defparam \Selector26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N8
cycloneive_lcell_comb \ShiftRight0~119 (
// Equation(s):
// \ShiftRight0~119_combout  = (Mux302 & ((Mux312 & ((\portB~49_combout ))) # (!Mux312 & (\portB~51_combout ))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB24),
	.datad(portB23),
	.cin(gnd),
	.combout(\ShiftRight0~119_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~119 .lut_mask = 16'hC840;
defparam \ShiftRight0~119 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N22
cycloneive_lcell_comb \ShiftRight0~120 (
// Equation(s):
// \ShiftRight0~120_combout  = (\ShiftRight0~119_combout ) # ((\ShiftRight0~55_combout  & !Mux302))

	.dataa(gnd),
	.datab(\ShiftRight0~55_combout ),
	.datac(Mux302),
	.datad(\ShiftRight0~119_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~120_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~120 .lut_mask = 16'hFF0C;
defparam \ShiftRight0~120 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N24
cycloneive_lcell_comb \ShiftRight0~117 (
// Equation(s):
// \ShiftRight0~117_combout  = (Mux312 & (((\portB~41_combout )) # (!Mux302))) # (!Mux312 & (Mux302 & (\portB~43_combout )))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB20),
	.datad(portB19),
	.cin(gnd),
	.combout(\ShiftRight0~117_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~117 .lut_mask = 16'hEA62;
defparam \ShiftRight0~117 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N2
cycloneive_lcell_comb \ShiftRight0~118 (
// Equation(s):
// \ShiftRight0~118_combout  = (Mux302 & (((\ShiftRight0~117_combout )))) # (!Mux302 & ((\ShiftRight0~117_combout  & (\portB~45_combout )) # (!\ShiftRight0~117_combout  & ((\portB~47_combout )))))

	.dataa(portB21),
	.datab(Mux302),
	.datac(portB22),
	.datad(\ShiftRight0~117_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~118_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~118 .lut_mask = 16'hEE30;
defparam \ShiftRight0~118 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N16
cycloneive_lcell_comb \Selector26~5 (
// Equation(s):
// \Selector26~5_combout  = (\Selector7~18_combout  & (\Selector7~10_combout )) # (!\Selector7~18_combout  & ((\Selector7~10_combout  & ((\ShiftRight0~118_combout ))) # (!\Selector7~10_combout  & (\ShiftRight0~120_combout ))))

	.dataa(\Selector7~18_combout ),
	.datab(\Selector7~10_combout ),
	.datac(\ShiftRight0~120_combout ),
	.datad(\ShiftRight0~118_combout ),
	.cin(gnd),
	.combout(\Selector26~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~5 .lut_mask = 16'hDC98;
defparam \Selector26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N6
cycloneive_lcell_comb \Selector26~6 (
// Equation(s):
// \Selector26~6_combout  = (\Selector7~18_combout  & ((\Selector26~5_combout  & ((\ShiftRight0~99_combout ))) # (!\Selector26~5_combout  & (\ShiftRight0~116_combout )))) # (!\Selector7~18_combout  & (\Selector26~5_combout ))

	.dataa(\Selector7~18_combout ),
	.datab(\Selector26~5_combout ),
	.datac(\ShiftRight0~116_combout ),
	.datad(\ShiftRight0~99_combout ),
	.cin(gnd),
	.combout(\Selector26~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~6 .lut_mask = 16'hEC64;
defparam \Selector26~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N16
cycloneive_lcell_comb \Selector19~0 (
// Equation(s):
// \Selector19~0_combout  = (\Selector0~35_combout  & ((Mux292 & (\ShiftRight0~29_combout )) # (!Mux292 & ((\ShiftRight0~33_combout )))))

	.dataa(Mux292),
	.datab(\Selector0~35_combout ),
	.datac(\ShiftRight0~29_combout ),
	.datad(\ShiftRight0~33_combout ),
	.cin(gnd),
	.combout(\Selector19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~0 .lut_mask = 16'hC480;
defparam \Selector19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N26
cycloneive_lcell_comb \Selector19~1 (
// Equation(s):
// \Selector19~1_combout  = (\Selector19~0_combout ) # ((\ShiftRight0~124_combout  & (\ShiftRight0~26_combout  & Selector22)))

	.dataa(\ShiftRight0~124_combout ),
	.datab(\ShiftRight0~26_combout ),
	.datac(Selector22),
	.datad(\Selector19~0_combout ),
	.cin(gnd),
	.combout(\Selector19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~1 .lut_mask = 16'hFF80;
defparam \Selector19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N10
cycloneive_lcell_comb \ShiftRight0~34 (
// Equation(s):
// \ShiftRight0~34_combout  = (!Mux302 & ((Mux312 & ((\portB~31_combout ))) # (!Mux312 & (\portB~33_combout ))))

	.dataa(Mux302),
	.datab(Mux312),
	.datac(portB15),
	.datad(portB14),
	.cin(gnd),
	.combout(\ShiftRight0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~34 .lut_mask = 16'h5410;
defparam \ShiftRight0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N8
cycloneive_lcell_comb \ShiftRight0~113 (
// Equation(s):
// \ShiftRight0~113_combout  = (Mux292 & ((\ShiftRight0~35_combout ) # ((\ShiftRight0~34_combout )))) # (!Mux292 & (((\ShiftRight0~46_combout ))))

	.dataa(\ShiftRight0~35_combout ),
	.datab(\ShiftRight0~34_combout ),
	.datac(Mux292),
	.datad(\ShiftRight0~46_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~113_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~113 .lut_mask = 16'hEFE0;
defparam \ShiftRight0~113 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N16
cycloneive_lcell_comb \Selector19~4 (
// Equation(s):
// \Selector19~4_combout  = (\portB~41_combout  & ((\Selector0~17_combout ) # ((Mux19 & \Selector0~18_combout ))))

	.dataa(portB19),
	.datab(\Selector0~17_combout ),
	.datac(Mux19),
	.datad(\Selector0~18_combout ),
	.cin(gnd),
	.combout(\Selector19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~4 .lut_mask = 16'hA888;
defparam \Selector19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N30
cycloneive_lcell_comb \Selector19~5 (
// Equation(s):
// \Selector19~5_combout  = (\Selector19~4_combout ) # ((!\portB~41_combout  & (!Mux19 & \Selector0~27_combout )))

	.dataa(portB19),
	.datab(\Selector19~4_combout ),
	.datac(Mux19),
	.datad(\Selector0~27_combout ),
	.cin(gnd),
	.combout(\Selector19~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~5 .lut_mask = 16'hCDCC;
defparam \Selector19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N20
cycloneive_lcell_comb \Selector19~6 (
// Equation(s):
// \Selector19~6_combout  = (\Selector19~5_combout ) # ((\Selector0~15_combout  & (\portB~41_combout  $ (Mux19))))

	.dataa(portB19),
	.datab(Mux19),
	.datac(\Selector19~5_combout ),
	.datad(\Selector0~15_combout ),
	.cin(gnd),
	.combout(\Selector19~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~6 .lut_mask = 16'hF6F0;
defparam \Selector19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N6
cycloneive_lcell_comb \Selector19~2 (
// Equation(s):
// \Selector19~2_combout  = (\Selector0~31_combout  & ((\Add0~24_combout ) # ((\Selector0~14_combout  & \Add1~24_combout )))) # (!\Selector0~31_combout  & (\Selector0~14_combout  & (\Add1~24_combout )))

	.dataa(\Selector0~31_combout ),
	.datab(\Selector0~14_combout ),
	.datac(\Add1~24_combout ),
	.datad(\Add0~24_combout ),
	.cin(gnd),
	.combout(\Selector19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~2 .lut_mask = 16'hEAC0;
defparam \Selector19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N28
cycloneive_lcell_comb \Selector19~3 (
// Equation(s):
// \Selector19~3_combout  = (\Selector19~2_combout ) # ((Mux19 & \Selector0~17_combout ))

	.dataa(gnd),
	.datab(Mux19),
	.datac(\Selector0~17_combout ),
	.datad(\Selector19~2_combout ),
	.cin(gnd),
	.combout(\Selector19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~3 .lut_mask = 16'hFFC0;
defparam \Selector19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N18
cycloneive_lcell_comb \Selector19~7 (
// Equation(s):
// \Selector19~7_combout  = (\Selector19~6_combout ) # ((\Selector19~3_combout ) # ((\ShiftRight0~113_combout  & \Selector16~9_combout )))

	.dataa(\ShiftRight0~113_combout ),
	.datab(\Selector19~6_combout ),
	.datac(\Selector16~9_combout ),
	.datad(\Selector19~3_combout ),
	.cin(gnd),
	.combout(\Selector19~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~7 .lut_mask = 16'hFFEC;
defparam \Selector19~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N2
cycloneive_lcell_comb \Selector20~1 (
// Equation(s):
// \Selector20~1_combout  = (cuifALUOP_0 & (!Mux28 & (\Selector1~8_combout  & Mux272)))

	.dataa(cuifALUOP_0),
	.datab(Mux28),
	.datac(\Selector1~8_combout ),
	.datad(Mux272),
	.cin(gnd),
	.combout(\Selector20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~1 .lut_mask = 16'h2000;
defparam \Selector20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N26
cycloneive_lcell_comb \Selector20~3 (
// Equation(s):
// \Selector20~3_combout  = (\Add0~22_combout  & ((\Selector0~31_combout ) # ((\Selector0~14_combout  & \Add1~22_combout )))) # (!\Add0~22_combout  & (((\Selector0~14_combout  & \Add1~22_combout ))))

	.dataa(\Add0~22_combout ),
	.datab(\Selector0~31_combout ),
	.datac(\Selector0~14_combout ),
	.datad(\Add1~22_combout ),
	.cin(gnd),
	.combout(\Selector20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~3 .lut_mask = 16'hF888;
defparam \Selector20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N18
cycloneive_lcell_comb \Selector20~4 (
// Equation(s):
// \Selector20~4_combout  = (\portB~43_combout  & ((\Selector0~17_combout ) # ((Mux20 & \Selector0~18_combout ))))

	.dataa(portB20),
	.datab(Mux20),
	.datac(\Selector0~18_combout ),
	.datad(\Selector0~17_combout ),
	.cin(gnd),
	.combout(\Selector20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~4 .lut_mask = 16'hAA80;
defparam \Selector20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N20
cycloneive_lcell_comb \Selector20~5 (
// Equation(s):
// \Selector20~5_combout  = (\Selector20~4_combout ) # ((\Selector0~27_combout  & (!Mux20 & !\portB~43_combout )))

	.dataa(\Selector0~27_combout ),
	.datab(Mux20),
	.datac(portB20),
	.datad(\Selector20~4_combout ),
	.cin(gnd),
	.combout(\Selector20~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~5 .lut_mask = 16'hFF02;
defparam \Selector20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N30
cycloneive_lcell_comb \Selector20~6 (
// Equation(s):
// \Selector20~6_combout  = (\Selector20~5_combout ) # ((\Selector0~15_combout  & (Mux20 $ (\portB~43_combout ))))

	.dataa(Mux20),
	.datab(portB20),
	.datac(\Selector0~15_combout ),
	.datad(\Selector20~5_combout ),
	.cin(gnd),
	.combout(\Selector20~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~6 .lut_mask = 16'hFF60;
defparam \Selector20~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N26
cycloneive_lcell_comb \Selector21~3 (
// Equation(s):
// \Selector21~3_combout  = (\portB~45_combout  & ((\Selector0~17_combout ) # ((Mux21 & \Selector0~18_combout ))))

	.dataa(Mux21),
	.datab(portB21),
	.datac(\Selector0~18_combout ),
	.datad(\Selector0~17_combout ),
	.cin(gnd),
	.combout(\Selector21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~3 .lut_mask = 16'hCC80;
defparam \Selector21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N0
cycloneive_lcell_comb \Selector21~4 (
// Equation(s):
// \Selector21~4_combout  = (\Selector21~3_combout ) # ((!Mux21 & (!\portB~45_combout  & \Selector0~27_combout )))

	.dataa(Mux21),
	.datab(portB21),
	.datac(\Selector21~3_combout ),
	.datad(\Selector0~27_combout ),
	.cin(gnd),
	.combout(\Selector21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~4 .lut_mask = 16'hF1F0;
defparam \Selector21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N6
cycloneive_lcell_comb \Selector21~5 (
// Equation(s):
// \Selector21~5_combout  = (\Selector21~4_combout ) # ((\Selector0~15_combout  & (Mux21 $ (\portB~45_combout ))))

	.dataa(Mux21),
	.datab(\Selector21~4_combout ),
	.datac(portB21),
	.datad(\Selector0~15_combout ),
	.cin(gnd),
	.combout(\Selector21~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~5 .lut_mask = 16'hDECC;
defparam \Selector21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N16
cycloneive_lcell_comb \Selector21~2 (
// Equation(s):
// \Selector21~2_combout  = (\Selector0~14_combout  & ((\Add1~20_combout ) # ((\Selector0~31_combout  & \Add0~20_combout )))) # (!\Selector0~14_combout  & (\Selector0~31_combout  & ((\Add0~20_combout ))))

	.dataa(\Selector0~14_combout ),
	.datab(\Selector0~31_combout ),
	.datac(\Add1~20_combout ),
	.datad(\Add0~20_combout ),
	.cin(gnd),
	.combout(\Selector21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~2 .lut_mask = 16'hECA0;
defparam \Selector21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N6
cycloneive_lcell_comb \Selector8~5 (
// Equation(s):
// \Selector8~5_combout  = (\portB~19_combout  & ((\Selector0~17_combout ) # ((Mux8 & \Selector0~18_combout ))))

	.dataa(Mux8),
	.datab(\Selector0~17_combout ),
	.datac(portB8),
	.datad(\Selector0~18_combout ),
	.cin(gnd),
	.combout(\Selector8~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~5 .lut_mask = 16'hE0C0;
defparam \Selector8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N28
cycloneive_lcell_comb \Selector8~6 (
// Equation(s):
// \Selector8~6_combout  = (\Selector8~5_combout ) # ((!Mux8 & (\Selector0~27_combout  & !\portB~19_combout )))

	.dataa(Mux8),
	.datab(\Selector0~27_combout ),
	.datac(portB8),
	.datad(\Selector8~5_combout ),
	.cin(gnd),
	.combout(\Selector8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~6 .lut_mask = 16'hFF04;
defparam \Selector8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N26
cycloneive_lcell_comb \Selector8~7 (
// Equation(s):
// \Selector8~7_combout  = (\Selector8~6_combout ) # ((\Selector0~15_combout  & (Mux8 $ (\portB~19_combout ))))

	.dataa(Mux8),
	.datab(\Selector0~15_combout ),
	.datac(portB8),
	.datad(\Selector8~6_combout ),
	.cin(gnd),
	.combout(\Selector8~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~7 .lut_mask = 16'hFF48;
defparam \Selector8~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N10
cycloneive_lcell_comb \Selector8~4 (
// Equation(s):
// \Selector8~4_combout  = (\Selector0~14_combout  & ((\Add1~46_combout ) # ((\Selector0~31_combout  & \Add0~46_combout )))) # (!\Selector0~14_combout  & (\Selector0~31_combout  & ((\Add0~46_combout ))))

	.dataa(\Selector0~14_combout ),
	.datab(\Selector0~31_combout ),
	.datac(\Add1~46_combout ),
	.datad(\Add0~46_combout ),
	.cin(gnd),
	.combout(\Selector8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~4 .lut_mask = 16'hECA0;
defparam \Selector8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N6
cycloneive_lcell_comb \Selector9~3 (
// Equation(s):
// \Selector9~3_combout  = (\portB~21_combout  & ((\Selector0~17_combout ) # ((Mux9 & \Selector0~18_combout ))))

	.dataa(Mux9),
	.datab(\Selector0~17_combout ),
	.datac(\Selector0~18_combout ),
	.datad(portB9),
	.cin(gnd),
	.combout(\Selector9~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~3 .lut_mask = 16'hEC00;
defparam \Selector9~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N24
cycloneive_lcell_comb \Selector9~4 (
// Equation(s):
// \Selector9~4_combout  = (\Selector9~3_combout ) # ((!Mux9 & (!\portB~21_combout  & \Selector0~27_combout )))

	.dataa(Mux9),
	.datab(portB9),
	.datac(\Selector0~27_combout ),
	.datad(\Selector9~3_combout ),
	.cin(gnd),
	.combout(\Selector9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~4 .lut_mask = 16'hFF10;
defparam \Selector9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N26
cycloneive_lcell_comb \Selector9~5 (
// Equation(s):
// \Selector9~5_combout  = (\Selector9~4_combout ) # ((\Selector0~15_combout  & (\portB~21_combout  $ (Mux9))))

	.dataa(portB9),
	.datab(\Selector0~15_combout ),
	.datac(Mux9),
	.datad(\Selector9~4_combout ),
	.cin(gnd),
	.combout(\Selector9~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~5 .lut_mask = 16'hFF48;
defparam \Selector9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N14
cycloneive_lcell_comb \Selector9~2 (
// Equation(s):
// \Selector9~2_combout  = (\Selector0~31_combout  & ((\Add0~44_combout ) # ((\Add1~44_combout  & \Selector0~14_combout )))) # (!\Selector0~31_combout  & (\Add1~44_combout  & ((\Selector0~14_combout ))))

	.dataa(\Selector0~31_combout ),
	.datab(\Add1~44_combout ),
	.datac(\Add0~44_combout ),
	.datad(\Selector0~14_combout ),
	.cin(gnd),
	.combout(\Selector9~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~2 .lut_mask = 16'hECA0;
defparam \Selector9~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N26
cycloneive_lcell_comb \Selector1~26 (
// Equation(s):
// \Selector1~26_combout  = (Mux292 & ((\ShiftLeft0~83_combout ) # ((\ShiftLeft0~82_combout )))) # (!Mux292 & (((\ShiftLeft0~87_combout ))))

	.dataa(Mux292),
	.datab(\ShiftLeft0~83_combout ),
	.datac(\ShiftLeft0~87_combout ),
	.datad(\ShiftLeft0~82_combout ),
	.cin(gnd),
	.combout(\Selector1~26_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~26 .lut_mask = 16'hFAD8;
defparam \Selector1~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N20
cycloneive_lcell_comb \Selector22~2 (
// Equation(s):
// \Selector22~2_combout  = (\Selector22~1_combout  & ((\Selector0~35_combout ) # ((\Selector20~1_combout  & \ShiftRight0~109_combout )))) # (!\Selector22~1_combout  & (\Selector20~1_combout  & (\ShiftRight0~109_combout )))

	.dataa(\Selector22~1_combout ),
	.datab(\Selector20~1_combout ),
	.datac(\ShiftRight0~109_combout ),
	.datad(\Selector0~35_combout ),
	.cin(gnd),
	.combout(\Selector22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~2 .lut_mask = 16'hEAC0;
defparam \Selector22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N24
cycloneive_lcell_comb \Selector22~5 (
// Equation(s):
// \Selector22~5_combout  = (\portB~47_combout  & ((\Selector0~17_combout ) # ((\Selector0~18_combout  & Mux22))))

	.dataa(\Selector0~18_combout ),
	.datab(Mux22),
	.datac(portB22),
	.datad(\Selector0~17_combout ),
	.cin(gnd),
	.combout(\Selector22~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~5 .lut_mask = 16'hF080;
defparam \Selector22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N22
cycloneive_lcell_comb \Selector22~6 (
// Equation(s):
// \Selector22~6_combout  = (\Selector22~5_combout ) # ((\Selector0~27_combout  & (!Mux22 & !\portB~47_combout )))

	.dataa(\Selector0~27_combout ),
	.datab(Mux22),
	.datac(portB22),
	.datad(\Selector22~5_combout ),
	.cin(gnd),
	.combout(\Selector22~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~6 .lut_mask = 16'hFF02;
defparam \Selector22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N12
cycloneive_lcell_comb \Selector22~7 (
// Equation(s):
// \Selector22~7_combout  = (\Selector22~6_combout ) # ((\Selector0~15_combout  & (Mux22 $ (\portB~47_combout ))))

	.dataa(\Selector22~6_combout ),
	.datab(Mux22),
	.datac(portB22),
	.datad(\Selector0~15_combout ),
	.cin(gnd),
	.combout(\Selector22~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~7 .lut_mask = 16'hBEAA;
defparam \Selector22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N16
cycloneive_lcell_comb \Selector22~3 (
// Equation(s):
// \Selector22~3_combout  = (\Selector0~14_combout  & ((\Add1~18_combout ) # ((\Selector0~31_combout  & \Add0~18_combout )))) # (!\Selector0~14_combout  & (\Selector0~31_combout  & ((\Add0~18_combout ))))

	.dataa(\Selector0~14_combout ),
	.datab(\Selector0~31_combout ),
	.datac(\Add1~18_combout ),
	.datad(\Add0~18_combout ),
	.cin(gnd),
	.combout(\Selector22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~3 .lut_mask = 16'hECA0;
defparam \Selector22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N2
cycloneive_lcell_comb \Selector22~4 (
// Equation(s):
// \Selector22~4_combout  = (\Selector22~3_combout ) # ((\Selector0~17_combout  & Mux22))

	.dataa(\Selector0~17_combout ),
	.datab(gnd),
	.datac(Mux22),
	.datad(\Selector22~3_combout ),
	.cin(gnd),
	.combout(\Selector22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~4 .lut_mask = 16'hFFA0;
defparam \Selector22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N28
cycloneive_lcell_comb \Selector30~2 (
// Equation(s):
// \Selector30~2_combout  = (Mux292 & ((\ShiftRight0~114_combout ) # ((\ShiftRight0~115_combout )))) # (!Mux292 & (((\ShiftRight0~118_combout ))))

	.dataa(\ShiftRight0~114_combout ),
	.datab(\ShiftRight0~115_combout ),
	.datac(Mux292),
	.datad(\ShiftRight0~118_combout ),
	.cin(gnd),
	.combout(\Selector30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~2 .lut_mask = 16'hEFE0;
defparam \Selector30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N20
cycloneive_lcell_comb \Selector22~8 (
// Equation(s):
// \Selector22~8_combout  = (\Selector30~2_combout  & ((\Selector16~9_combout ) # ((\Selector16~1_combout  & \ShiftLeft0~100_combout )))) # (!\Selector30~2_combout  & (\Selector16~1_combout  & ((\ShiftLeft0~100_combout ))))

	.dataa(\Selector30~2_combout ),
	.datab(\Selector16~1_combout ),
	.datac(\Selector16~9_combout ),
	.datad(\ShiftLeft0~100_combout ),
	.cin(gnd),
	.combout(\Selector22~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~8 .lut_mask = 16'hECA0;
defparam \Selector22~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N22
cycloneive_lcell_comb \Selector30~8 (
// Equation(s):
// \Selector30~8_combout  = (\Selector0~5_combout ) # ((\portB~63_combout  & (\Selector0~6_combout )) # (!\portB~63_combout  & ((\Selector0~11_combout ))))

	.dataa(\Selector0~6_combout ),
	.datab(\Selector0~11_combout ),
	.datac(\Selector0~5_combout ),
	.datad(portB30),
	.cin(gnd),
	.combout(\Selector30~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~8 .lut_mask = 16'hFAFC;
defparam \Selector30~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N20
cycloneive_lcell_comb \Selector30~3 (
// Equation(s):
// \Selector30~3_combout  = (\portB~63_combout  & ((\Selector0~5_combout ) # ((!Mux302 & \Selector0~11_combout ))))

	.dataa(portB30),
	.datab(Mux302),
	.datac(\Selector0~5_combout ),
	.datad(\Selector0~11_combout ),
	.cin(gnd),
	.combout(\Selector30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~3 .lut_mask = 16'hA2A0;
defparam \Selector30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N10
cycloneive_lcell_comb \Selector30~4 (
// Equation(s):
// \Selector30~4_combout  = (\Selector4~0_combout  & (!Mux272 & (\Selector1~20_combout  & \ShiftLeft0~19_combout )))

	.dataa(\Selector4~0_combout ),
	.datab(Mux272),
	.datac(\Selector1~20_combout ),
	.datad(\ShiftLeft0~19_combout ),
	.cin(gnd),
	.combout(\Selector30~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~4 .lut_mask = 16'h2000;
defparam \Selector30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N12
cycloneive_lcell_comb \Selector30~5 (
// Equation(s):
// \Selector30~5_combout  = (\Add0~2_combout  & ((\Selector0~10_combout ) # ((\Selector0~8_combout  & \Add1~2_combout )))) # (!\Add0~2_combout  & (\Selector0~8_combout  & ((\Add1~2_combout ))))

	.dataa(\Add0~2_combout ),
	.datab(\Selector0~8_combout ),
	.datac(\Selector0~10_combout ),
	.datad(\Add1~2_combout ),
	.cin(gnd),
	.combout(\Selector30~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~5 .lut_mask = 16'hECA0;
defparam \Selector30~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N18
cycloneive_lcell_comb \Selector30~6 (
// Equation(s):
// \Selector30~6_combout  = (\Selector30~5_combout ) # ((!\portB~63_combout  & (!Mux302 & \Selector0~7_combout )))

	.dataa(portB30),
	.datab(Mux302),
	.datac(\Selector0~7_combout ),
	.datad(\Selector30~5_combout ),
	.cin(gnd),
	.combout(\Selector30~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~6 .lut_mask = 16'hFF10;
defparam \Selector30~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N4
cycloneive_lcell_comb \Selector30~7 (
// Equation(s):
// \Selector30~7_combout  = (\Selector30~3_combout ) # ((\Selector30~4_combout ) # (\Selector30~6_combout ))

	.dataa(gnd),
	.datab(\Selector30~3_combout ),
	.datac(\Selector30~4_combout ),
	.datad(\Selector30~6_combout ),
	.cin(gnd),
	.combout(\Selector30~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~7 .lut_mask = 16'hFFFC;
defparam \Selector30~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N14
cycloneive_lcell_comb \Selector30~15 (
// Equation(s):
// \Selector30~15_combout  = (Mux272 & (\Selector0~13_combout  & (\ShiftRight0~112_combout  & !\ShiftRight0~22_combout )))

	.dataa(Mux272),
	.datab(\Selector0~13_combout ),
	.datac(\ShiftRight0~112_combout ),
	.datad(\ShiftRight0~22_combout ),
	.cin(gnd),
	.combout(\Selector30~15_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~15 .lut_mask = 16'h0080;
defparam \Selector30~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N8
cycloneive_lcell_comb \Selector30~9 (
// Equation(s):
// \Selector30~9_combout  = (\Selector30~7_combout ) # ((\Selector30~15_combout ) # ((\Selector30~8_combout  & Mux302)))

	.dataa(\Selector30~8_combout ),
	.datab(Mux302),
	.datac(\Selector30~7_combout ),
	.datad(\Selector30~15_combout ),
	.cin(gnd),
	.combout(\Selector30~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~9 .lut_mask = 16'hFFF8;
defparam \Selector30~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N2
cycloneive_lcell_comb \Selector30~11 (
// Equation(s):
// \Selector30~11_combout  = (!Mux302 & ((Mux312 & ((\portB~61_combout ))) # (!Mux312 & (\portB~63_combout ))))

	.dataa(Mux312),
	.datab(Mux302),
	.datac(portB30),
	.datad(portB29),
	.cin(gnd),
	.combout(\Selector30~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~11 .lut_mask = 16'h3210;
defparam \Selector30~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N12
cycloneive_lcell_comb \Selector30~12 (
// Equation(s):
// \Selector30~12_combout  = (!Mux292 & ((\Selector30~11_combout ) # ((\ShiftRight0~59_combout  & Mux302))))

	.dataa(\ShiftRight0~59_combout ),
	.datab(Mux302),
	.datac(\Selector30~11_combout ),
	.datad(Mux292),
	.cin(gnd),
	.combout(\Selector30~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~12 .lut_mask = 16'h00F8;
defparam \Selector30~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N26
cycloneive_lcell_comb \Selector30~10 (
// Equation(s):
// \Selector30~10_combout  = (Mux292 & ((\ShiftRight0~119_combout ) # ((\ShiftRight0~55_combout  & !Mux302))))

	.dataa(Mux292),
	.datab(\ShiftRight0~55_combout ),
	.datac(Mux302),
	.datad(\ShiftRight0~119_combout ),
	.cin(gnd),
	.combout(\Selector30~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~10 .lut_mask = 16'hAA08;
defparam \Selector30~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N10
cycloneive_lcell_comb \Selector30~13 (
// Equation(s):
// \Selector30~13_combout  = (Mux28 & (((\Selector30~2_combout )))) # (!Mux28 & ((\Selector30~12_combout ) # ((\Selector30~10_combout ))))

	.dataa(\Selector30~12_combout ),
	.datab(Mux28),
	.datac(\Selector30~10_combout ),
	.datad(\Selector30~2_combout ),
	.cin(gnd),
	.combout(\Selector30~13_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~13 .lut_mask = 16'hFE32;
defparam \Selector30~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N6
cycloneive_lcell_comb \ShiftRight0~121 (
// Equation(s):
// \ShiftRight0~121_combout  = (Mux292 & (\ShiftRight0~46_combout )) # (!Mux292 & ((\ShiftRight0~48_combout )))

	.dataa(gnd),
	.datab(Mux292),
	.datac(\ShiftRight0~46_combout ),
	.datad(\ShiftRight0~48_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~121_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~121 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~121 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N8
cycloneive_lcell_comb \Selector23~6 (
// Equation(s):
// \Selector23~6_combout  = (\portB~49_combout  & ((\Selector0~17_combout ) # ((\Selector0~18_combout  & Mux23))))

	.dataa(\Selector0~17_combout ),
	.datab(portB23),
	.datac(\Selector0~18_combout ),
	.datad(Mux23),
	.cin(gnd),
	.combout(\Selector23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~6 .lut_mask = 16'hC888;
defparam \Selector23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N30
cycloneive_lcell_comb \Selector23~7 (
// Equation(s):
// \Selector23~7_combout  = (\Selector23~6_combout ) # ((\Selector0~27_combout  & (!\portB~49_combout  & !Mux23)))

	.dataa(\Selector0~27_combout ),
	.datab(portB23),
	.datac(\Selector23~6_combout ),
	.datad(Mux23),
	.cin(gnd),
	.combout(\Selector23~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~7 .lut_mask = 16'hF0F2;
defparam \Selector23~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N4
cycloneive_lcell_comb \Selector23~8 (
// Equation(s):
// \Selector23~8_combout  = (\Selector23~7_combout ) # ((\Selector0~15_combout  & (Mux23 $ (\portB~49_combout ))))

	.dataa(Mux23),
	.datab(portB23),
	.datac(\Selector23~7_combout ),
	.datad(\Selector0~15_combout ),
	.cin(gnd),
	.combout(\Selector23~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~8 .lut_mask = 16'hF6F0;
defparam \Selector23~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N10
cycloneive_lcell_comb \Selector23~5 (
// Equation(s):
// \Selector23~5_combout  = (\Selector0~14_combout  & ((\Add1~16_combout ) # ((\Add0~16_combout  & \Selector0~31_combout )))) # (!\Selector0~14_combout  & (\Add0~16_combout  & (\Selector0~31_combout )))

	.dataa(\Selector0~14_combout ),
	.datab(\Add0~16_combout ),
	.datac(\Selector0~31_combout ),
	.datad(\Add1~16_combout ),
	.cin(gnd),
	.combout(\Selector23~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~5 .lut_mask = 16'hEAC0;
defparam \Selector23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N14
cycloneive_lcell_comb \Selector23~9 (
// Equation(s):
// \Selector23~9_combout  = (\Selector23~8_combout ) # ((\Selector23~5_combout ) # ((\Selector0~17_combout  & Mux23)))

	.dataa(\Selector0~17_combout ),
	.datab(Mux23),
	.datac(\Selector23~8_combout ),
	.datad(\Selector23~5_combout ),
	.cin(gnd),
	.combout(\Selector23~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~9 .lut_mask = 16'hFFF8;
defparam \Selector23~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N20
cycloneive_lcell_comb \Equal0~2 (
// Equation(s):
// \Equal0~2_combout  = (!Selector41 & (!Selector2 & !Selector1))

	.dataa(Selector41),
	.datab(gnd),
	.datac(Selector2),
	.datad(Selector1),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~2 .lut_mask = 16'h0005;
defparam \Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N26
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (!Selector15 & (!Selector103 & (!Selector28 & !Selector291)))

	.dataa(Selector15),
	.datab(Selector103),
	.datac(Selector28),
	.datad(Selector291),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h0001;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N0
cycloneive_lcell_comb \Equal0~1 (
// Equation(s):
// \Equal0~1_combout  = (!Selector7 & (!Selector3 & (\Equal0~0_combout  & !Selector111)))

	.dataa(Selector7),
	.datab(Selector3),
	.datac(\Equal0~0_combout ),
	.datad(Selector111),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~1 .lut_mask = 16'h0010;
defparam \Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N22
cycloneive_lcell_comb \Equal0~3 (
// Equation(s):
// \Equal0~3_combout  = (!Selector311 & (!Selector0 & (\Equal0~2_combout  & \Equal0~1_combout )))

	.dataa(Selector311),
	.datab(Selector0),
	.datac(\Equal0~2_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~3 .lut_mask = 16'h1000;
defparam \Equal0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N30
cycloneive_lcell_comb \Equal0~10 (
// Equation(s):
// \Equal0~10_combout  = (!Selector232 & (!Selector231 & (!Selector23 & !Selector30)))

	.dataa(Selector232),
	.datab(Selector231),
	.datac(Selector23),
	.datad(Selector30),
	.cin(gnd),
	.combout(\Equal0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~10 .lut_mask = 16'h0001;
defparam \Equal0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N20
cycloneive_lcell_comb \Equal0~5 (
// Equation(s):
// \Equal0~5_combout  = (!Selector16 & (!Selector27 & (!Selector143 & !Selector25)))

	.dataa(Selector16),
	.datab(Selector27),
	.datac(Selector143),
	.datad(Selector25),
	.cin(gnd),
	.combout(\Equal0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~5 .lut_mask = 16'h0001;
defparam \Equal0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N0
cycloneive_lcell_comb \Equal0~7 (
// Equation(s):
// \Equal0~7_combout  = (!Selector202 & (!Selector20 & (!Selector19 & !Selector201)))

	.dataa(Selector202),
	.datab(Selector20),
	.datac(Selector19),
	.datad(Selector201),
	.cin(gnd),
	.combout(\Equal0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~7 .lut_mask = 16'h0001;
defparam \Equal0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N4
cycloneive_lcell_comb \Equal0~4 (
// Equation(s):
// \Equal0~4_combout  = (!Selector12 & (!Selector13 & (!Selector242 & !Selector51)))

	.dataa(Selector12),
	.datab(Selector13),
	.datac(Selector242),
	.datad(Selector51),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~4 .lut_mask = 16'h0001;
defparam \Equal0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N2
cycloneive_lcell_comb \Equal0~6 (
// Equation(s):
// \Equal0~6_combout  = (!Selector17 & (!Selector6 & (!Selector18 & !Selector261)))

	.dataa(Selector17),
	.datab(Selector6),
	.datac(Selector18),
	.datad(Selector261),
	.cin(gnd),
	.combout(\Equal0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~6 .lut_mask = 16'h0001;
defparam \Equal0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N8
cycloneive_lcell_comb \Equal0~8 (
// Equation(s):
// \Equal0~8_combout  = (\Equal0~5_combout  & (\Equal0~7_combout  & (\Equal0~4_combout  & \Equal0~6_combout )))

	.dataa(\Equal0~5_combout ),
	.datab(\Equal0~7_combout ),
	.datac(\Equal0~4_combout ),
	.datad(\Equal0~6_combout ),
	.cin(gnd),
	.combout(\Equal0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~8 .lut_mask = 16'h8000;
defparam \Equal0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N6
cycloneive_lcell_comb \Equal0~9 (
// Equation(s):
// \Equal0~9_combout  = (!Selector213 & (!Selector221 & (!Selector84 & !Selector93)))

	.dataa(Selector213),
	.datab(Selector221),
	.datac(Selector84),
	.datad(Selector93),
	.cin(gnd),
	.combout(\Equal0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~9 .lut_mask = 16'h0001;
defparam \Equal0~9 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module control_unit (
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	instr_30,
	ccifiwait_0,
	dcifimemload_30,
	instr_31,
	dcifimemload_31,
	instr_27,
	dcifimemload_27,
	instr_26,
	dcifimemload_26,
	instr_29,
	dcifimemload_29,
	instr_28,
	dcifimemload_28,
	Equal6,
	Equal0,
	dcifimemload_3,
	dcifimemload_4,
	dcifimemload_2,
	dcifimemload_5,
	dcifimemload_0,
	dcifimemload_1,
	always0,
	cuifRegWEN,
	Equal7,
	Equal3,
	cuifALUOP_3,
	cuifALUOP_2,
	cuifALUOP_1,
	cuifALUOP_0,
	Equal01,
	Equal2,
	Equal31,
	cuifPCSrc_0,
	dcifdhit,
	cuifPCSrc_1,
	cuifMemtoReg_0,
	cuifMemtoReg_1,
	cuifRegWEN1,
	cuifALUOP_21,
	devpor,
	devclrn,
	devoe);
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	instr_30;
input 	ccifiwait_0;
input 	dcifimemload_30;
input 	instr_31;
input 	dcifimemload_31;
input 	instr_27;
input 	dcifimemload_27;
input 	instr_26;
input 	dcifimemload_26;
input 	instr_29;
input 	dcifimemload_29;
input 	instr_28;
input 	dcifimemload_28;
output 	Equal6;
output 	Equal0;
input 	dcifimemload_3;
input 	dcifimemload_4;
input 	dcifimemload_2;
input 	dcifimemload_5;
input 	dcifimemload_0;
input 	dcifimemload_1;
output 	always0;
output 	cuifRegWEN;
output 	Equal7;
output 	Equal3;
output 	cuifALUOP_3;
output 	cuifALUOP_2;
output 	cuifALUOP_1;
output 	cuifALUOP_0;
input 	Equal01;
output 	Equal2;
output 	Equal31;
output 	cuifPCSrc_0;
input 	dcifdhit;
output 	cuifPCSrc_1;
output 	cuifMemtoReg_0;
output 	cuifMemtoReg_1;
output 	cuifRegWEN1;
output 	cuifALUOP_21;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \always0~2_combout ;
wire \Equal6~0_combout ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal2~0_combout ;
wire \Equal2~1_combout ;
wire \always0~0_combout ;
wire \cuif.ALUOP[1]~2_combout ;
wire \cuif.ALUOP[1]~3_combout ;
wire \Equal26~0_combout ;
wire \Equal8~0_combout ;
wire \cuif.ALUOP[3]~4_combout ;
wire \Equal25~0_combout ;
wire \cuif.ALUOP[3]~7_combout ;
wire \cuif.ALUOP[3]~5_combout ;
wire \cuif.ALUOP[3]~6_combout ;
wire \cuif.ALUOP[2]~9_combout ;
wire \cuif.ALUOP[2]~10_combout ;
wire \cuif.ALUOP[1]~12_combout ;
wire \cuif.ALUOP[1]~13_combout ;
wire \cuif.ALUOP[1]~14_combout ;
wire \Equal11~2_combout ;
wire \cuif.ALUOP[1]~15_combout ;
wire \cuif.ALUOP[0]~21_combout ;
wire \cuif.ALUOP[0]~22_combout ;
wire \cuif.ALUOP[0]~18_combout ;
wire \Equal7~1_combout ;
wire \cuif.ALUOP[0]~17_combout ;
wire \Equal4~0_combout ;
wire \cuif.PCSrc[0]~0_combout ;
wire \Equal10~0_combout ;
wire \cuif.RegWEN~1_combout ;


// Location: LCCOMB_X57_Y29_N10
cycloneive_lcell_comb \always0~2 (
// Equation(s):
// \always0~2_combout  = (dcifimemload_31 & (dcifimemload_27 & (dcifimemload_26))) # (!dcifimemload_31 & (!dcifimemload_27 & ((dcifimemload_29))))

	.dataa(dcifimemload_31),
	.datab(dcifimemload_27),
	.datac(dcifimemload_26),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
// synopsys translate_off
defparam \always0~2 .lut_mask = 16'h9180;
defparam \always0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N22
cycloneive_lcell_comb \Equal6~1 (
// Equation(s):
// Equal6 = (dcifimemload_29 & (dcifimemload_28 & \Equal6~0_combout ))

	.dataa(gnd),
	.datab(dcifimemload_29),
	.datac(dcifimemload_28),
	.datad(\Equal6~0_combout ),
	.cin(gnd),
	.combout(Equal6),
	.cout());
// synopsys translate_off
defparam \Equal6~1 .lut_mask = 16'hC000;
defparam \Equal6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N30
cycloneive_lcell_comb \Equal0~2 (
// Equation(s):
// Equal0 = (\Equal0~1_combout  & (\Equal2~1_combout  & (!dcifimemload_29 & !dcifimemload_27)))

	.dataa(\Equal0~1_combout ),
	.datab(\Equal2~1_combout ),
	.datac(dcifimemload_29),
	.datad(dcifimemload_27),
	.cin(gnd),
	.combout(Equal0),
	.cout());
// synopsys translate_off
defparam \Equal0~2 .lut_mask = 16'h0008;
defparam \Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N24
cycloneive_lcell_comb \always0~1 (
// Equation(s):
// always0 = (!dcifimemload_5 & (!dcifimemload_0 & (!dcifimemload_1 & \always0~0_combout )))

	.dataa(dcifimemload_5),
	.datab(dcifimemload_0),
	.datac(dcifimemload_1),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(always0),
	.cout());
// synopsys translate_off
defparam \always0~1 .lut_mask = 16'h0100;
defparam \always0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N0
cycloneive_lcell_comb \cuif.RegWEN~0 (
// Equation(s):
// cuifRegWEN = ((!\cuif.ALUOP[1]~3_combout ) # (!dcifimemload_28)) # (!\Equal0~1_combout )

	.dataa(gnd),
	.datab(\Equal0~1_combout ),
	.datac(dcifimemload_28),
	.datad(\cuif.ALUOP[1]~3_combout ),
	.cin(gnd),
	.combout(cuifRegWEN),
	.cout());
// synopsys translate_off
defparam \cuif.RegWEN~0 .lut_mask = 16'h3FFF;
defparam \cuif.RegWEN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N30
cycloneive_lcell_comb \Equal7~0 (
// Equation(s):
// Equal7 = (!dcifimemload_31 & (dcifimemload_29 & (!dcifimemload_30 & dcifimemload_28)))

	.dataa(dcifimemload_31),
	.datab(dcifimemload_29),
	.datac(dcifimemload_30),
	.datad(dcifimemload_28),
	.cin(gnd),
	.combout(Equal7),
	.cout());
// synopsys translate_off
defparam \Equal7~0 .lut_mask = 16'h0400;
defparam \Equal7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N14
cycloneive_lcell_comb \Equal3~0 (
// Equation(s):
// Equal3 = (dcifimemload_26 & (!dcifimemload_30 & (dcifimemload_27 & !dcifimemload_28)))

	.dataa(dcifimemload_26),
	.datab(dcifimemload_30),
	.datac(dcifimemload_27),
	.datad(dcifimemload_28),
	.cin(gnd),
	.combout(Equal3),
	.cout());
// synopsys translate_off
defparam \Equal3~0 .lut_mask = 16'h0020;
defparam \Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N6
cycloneive_lcell_comb \cuif.ALUOP[3]~8 (
// Equation(s):
// cuifALUOP_3 = (\cuif.ALUOP[3]~5_combout ) # ((\cuif.ALUOP[3]~6_combout ) # ((\Equal26~0_combout  & \cuif.ALUOP[3]~7_combout )))

	.dataa(\Equal26~0_combout ),
	.datab(\cuif.ALUOP[3]~7_combout ),
	.datac(\cuif.ALUOP[3]~5_combout ),
	.datad(\cuif.ALUOP[3]~6_combout ),
	.cin(gnd),
	.combout(cuifALUOP_3),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[3]~8 .lut_mask = 16'hFFF8;
defparam \cuif.ALUOP[3]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N8
cycloneive_lcell_comb \cuif.ALUOP[2]~11 (
// Equation(s):
// cuifALUOP_2 = (\cuif.ALUOP[2]~10_combout ) # ((!\Equal26~0_combout  & \cuif.ALUOP[3]~7_combout ))

	.dataa(gnd),
	.datab(\Equal26~0_combout ),
	.datac(\cuif.ALUOP[2]~10_combout ),
	.datad(\cuif.ALUOP[3]~7_combout ),
	.cin(gnd),
	.combout(cuifALUOP_2),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[2]~11 .lut_mask = 16'hF3F0;
defparam \cuif.ALUOP[2]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N30
cycloneive_lcell_comb \cuif.ALUOP[1]~16 (
// Equation(s):
// cuifALUOP_1 = (\Equal11~2_combout ) # ((\Equal0~1_combout  & ((\cuif.ALUOP[1]~14_combout ) # (\cuif.ALUOP[1]~15_combout ))))

	.dataa(\cuif.ALUOP[1]~14_combout ),
	.datab(\Equal11~2_combout ),
	.datac(\Equal0~1_combout ),
	.datad(\cuif.ALUOP[1]~15_combout ),
	.cin(gnd),
	.combout(cuifALUOP_1),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[1]~16 .lut_mask = 16'hFCEC;
defparam \cuif.ALUOP[1]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N6
cycloneive_lcell_comb \cuif.ALUOP[0]~19 (
// Equation(s):
// cuifALUOP_0 = ((\Equal26~0_combout ) # ((\cuif.ALUOP[0]~18_combout ) # (\cuif.ALUOP[0]~17_combout ))) # (!cuifRegWEN)

	.dataa(cuifRegWEN),
	.datab(\Equal26~0_combout ),
	.datac(\cuif.ALUOP[0]~18_combout ),
	.datad(\cuif.ALUOP[0]~17_combout ),
	.cin(gnd),
	.combout(cuifALUOP_0),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[0]~19 .lut_mask = 16'hFFFD;
defparam \cuif.ALUOP[0]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N16
cycloneive_lcell_comb \Equal2~2 (
// Equation(s):
// Equal2 = (!dcifimemload_29 & (\Equal2~1_combout  & (\Equal0~1_combout  & dcifimemload_27)))

	.dataa(dcifimemload_29),
	.datab(\Equal2~1_combout ),
	.datac(\Equal0~1_combout ),
	.datad(dcifimemload_27),
	.cin(gnd),
	.combout(Equal2),
	.cout());
// synopsys translate_off
defparam \Equal2~2 .lut_mask = 16'h4000;
defparam \Equal2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N16
cycloneive_lcell_comb \Equal3~1 (
// Equation(s):
// Equal31 = (!dcifimemload_31 & (Equal3 & !dcifimemload_29))

	.dataa(dcifimemload_31),
	.datab(gnd),
	.datac(Equal3),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(Equal31),
	.cout());
// synopsys translate_off
defparam \Equal3~1 .lut_mask = 16'h0050;
defparam \Equal3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N30
cycloneive_lcell_comb \cuif.PCSrc[0]~1 (
// Equation(s):
// cuifPCSrc_0 = (!always0 & ((dcifimemload_26 $ (!Equal0)) # (!\cuif.PCSrc[0]~0_combout )))

	.dataa(dcifimemload_26),
	.datab(\cuif.PCSrc[0]~0_combout ),
	.datac(always0),
	.datad(Equal01),
	.cin(gnd),
	.combout(cuifPCSrc_0),
	.cout());
// synopsys translate_off
defparam \cuif.PCSrc[0]~1 .lut_mask = 16'h0B07;
defparam \cuif.PCSrc[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N18
cycloneive_lcell_comb \cuif.PCSrc[1]~2 (
// Equation(s):
// cuifPCSrc_1 = (Equal31) # ((always0) # (Equal2))

	.dataa(gnd),
	.datab(Equal31),
	.datac(always0),
	.datad(Equal2),
	.cin(gnd),
	.combout(cuifPCSrc_1),
	.cout());
// synopsys translate_off
defparam \cuif.PCSrc[1]~2 .lut_mask = 16'hFFFC;
defparam \cuif.PCSrc[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N16
cycloneive_lcell_comb \cuif.MemtoReg[0]~0 (
// Equation(s):
// cuifMemtoReg_0 = (\Equal11~2_combout  & (((Equal31 & !\Equal10~0_combout )) # (!dcifimemload_29))) # (!\Equal11~2_combout  & (((Equal31 & !\Equal10~0_combout ))))

	.dataa(\Equal11~2_combout ),
	.datab(dcifimemload_29),
	.datac(Equal31),
	.datad(\Equal10~0_combout ),
	.cin(gnd),
	.combout(cuifMemtoReg_0),
	.cout());
// synopsys translate_off
defparam \cuif.MemtoReg[0]~0 .lut_mask = 16'h22F2;
defparam \cuif.MemtoReg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N14
cycloneive_lcell_comb \cuif.MemtoReg[1]~1 (
// Equation(s):
// cuifMemtoReg_1 = (Equal31 & ((dcifimemload_29) # ((!\Equal11~2_combout )))) # (!Equal31 & (\Equal10~0_combout  & ((dcifimemload_29) # (!\Equal11~2_combout ))))

	.dataa(Equal31),
	.datab(dcifimemload_29),
	.datac(\Equal11~2_combout ),
	.datad(\Equal10~0_combout ),
	.cin(gnd),
	.combout(cuifMemtoReg_1),
	.cout());
// synopsys translate_off
defparam \cuif.MemtoReg[1]~1 .lut_mask = 16'hCF8A;
defparam \cuif.MemtoReg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N10
cycloneive_lcell_comb \cuif.RegWEN~2 (
// Equation(s):
// cuifRegWEN1 = (!Equal6 & (!Equal2 & (cuifRegWEN & \cuif.RegWEN~1_combout )))

	.dataa(Equal6),
	.datab(Equal2),
	.datac(cuifRegWEN),
	.datad(\cuif.RegWEN~1_combout ),
	.cin(gnd),
	.combout(cuifRegWEN1),
	.cout());
// synopsys translate_off
defparam \cuif.RegWEN~2 .lut_mask = 16'h1000;
defparam \cuif.RegWEN~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N14
cycloneive_lcell_comb \cuif.ALUOP[2]~20 (
// Equation(s):
// cuifALUOP_21 = (!Equal0 & (((!\cuif.ALUOP[1]~3_combout ) # (!\Equal0~1_combout )) # (!dcifimemload_28)))

	.dataa(dcifimemload_28),
	.datab(\Equal0~1_combout ),
	.datac(Equal0),
	.datad(\cuif.ALUOP[1]~3_combout ),
	.cin(gnd),
	.combout(cuifALUOP_21),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[2]~20 .lut_mask = 16'h070F;
defparam \cuif.ALUOP[2]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N20
cycloneive_lcell_comb \Equal6~0 (
// Equation(s):
// \Equal6~0_combout  = (dcifimemload_30 & (dcifimemload_31 & (dcifimemload_26 & dcifimemload_27)))

	.dataa(dcifimemload_30),
	.datab(dcifimemload_31),
	.datac(dcifimemload_26),
	.datad(dcifimemload_27),
	.cin(gnd),
	.combout(\Equal6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal6~0 .lut_mask = 16'h8000;
defparam \Equal6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N4
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (!instr_30 & !instr_31)

	.dataa(gnd),
	.datab(gnd),
	.datac(instr_30),
	.datad(instr_31),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h000F;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N28
cycloneive_lcell_comb \Equal0~1 (
// Equation(s):
// \Equal0~1_combout  = (ccifiwait_0 & (((!ramiframload_30 & !ramiframload_31)))) # (!ccifiwait_0 & (\Equal0~0_combout ))

	.dataa(\Equal0~0_combout ),
	.datab(ccifiwait_0),
	.datac(ramiframload_30),
	.datad(ramiframload_31),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~1 .lut_mask = 16'h222E;
defparam \Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N22
cycloneive_lcell_comb \Equal2~0 (
// Equation(s):
// \Equal2~0_combout  = (!instr_26 & !instr_28)

	.dataa(gnd),
	.datab(gnd),
	.datac(instr_26),
	.datad(instr_28),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~0 .lut_mask = 16'h000F;
defparam \Equal2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N16
cycloneive_lcell_comb \Equal2~1 (
// Equation(s):
// \Equal2~1_combout  = (ccifiwait_0 & (((!ramiframload_26 & !ramiframload_28)))) # (!ccifiwait_0 & (\Equal2~0_combout ))

	.dataa(\Equal2~0_combout ),
	.datab(ramiframload_26),
	.datac(ramiframload_28),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~1 .lut_mask = 16'h03AA;
defparam \Equal2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N28
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// \always0~0_combout  = (!dcifimemload_2 & (dcifimemload_3 & (!dcifimemload_4 & Equal0)))

	.dataa(dcifimemload_2),
	.datab(dcifimemload_3),
	.datac(dcifimemload_4),
	.datad(Equal0),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'h0400;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N18
cycloneive_lcell_comb \cuif.ALUOP[1]~2 (
// Equation(s):
// \cuif.ALUOP[1]~2_combout  = (!instr_27 & !instr_29)

	.dataa(gnd),
	.datab(gnd),
	.datac(instr_27),
	.datad(instr_29),
	.cin(gnd),
	.combout(\cuif.ALUOP[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[1]~2 .lut_mask = 16'h000F;
defparam \cuif.ALUOP[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N26
cycloneive_lcell_comb \cuif.ALUOP[1]~3 (
// Equation(s):
// \cuif.ALUOP[1]~3_combout  = (ccifiwait_0 & (!ramiframload_27 & ((!ramiframload_29)))) # (!ccifiwait_0 & (((\cuif.ALUOP[1]~2_combout ))))

	.dataa(ramiframload_27),
	.datab(\cuif.ALUOP[1]~2_combout ),
	.datac(ccifiwait_0),
	.datad(ramiframload_29),
	.cin(gnd),
	.combout(\cuif.ALUOP[1]~3_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[1]~3 .lut_mask = 16'h0C5C;
defparam \cuif.ALUOP[1]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N0
cycloneive_lcell_comb \Equal26~0 (
// Equation(s):
// \Equal26~0_combout  = (!dcifimemload_31 & (Equal3 & dcifimemload_29))

	.dataa(dcifimemload_31),
	.datab(gnd),
	.datac(Equal3),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(\Equal26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal26~0 .lut_mask = 16'h5000;
defparam \Equal26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N24
cycloneive_lcell_comb \Equal8~0 (
// Equation(s):
// \Equal8~0_combout  = (!dcifimemload_26 & (!dcifimemload_27 & Equal7))

	.dataa(dcifimemload_26),
	.datab(dcifimemload_27),
	.datac(Equal7),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal8~0 .lut_mask = 16'h1010;
defparam \Equal8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N2
cycloneive_lcell_comb \cuif.ALUOP[3]~4 (
// Equation(s):
// \cuif.ALUOP[3]~4_combout  = (!\Equal8~0_combout  & (((dcifimemload_30) # (dcifimemload_28)) # (!\always0~2_combout )))

	.dataa(\always0~2_combout ),
	.datab(dcifimemload_30),
	.datac(dcifimemload_28),
	.datad(\Equal8~0_combout ),
	.cin(gnd),
	.combout(\cuif.ALUOP[3]~4_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[3]~4 .lut_mask = 16'h00FD;
defparam \cuif.ALUOP[3]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N6
cycloneive_lcell_comb \Equal25~0 (
// Equation(s):
// \Equal25~0_combout  = (dcifimemload_29 & (\Equal2~1_combout  & (\Equal0~1_combout  & dcifimemload_27)))

	.dataa(dcifimemload_29),
	.datab(\Equal2~1_combout ),
	.datac(\Equal0~1_combout ),
	.datad(dcifimemload_27),
	.cin(gnd),
	.combout(\Equal25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal25~0 .lut_mask = 16'h8000;
defparam \Equal25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N16
cycloneive_lcell_comb \cuif.ALUOP[3]~7 (
// Equation(s):
// \cuif.ALUOP[3]~7_combout  = (cuifRegWEN & (\cuif.ALUOP[3]~4_combout  & (!\Equal25~0_combout  & !Equal0)))

	.dataa(cuifRegWEN),
	.datab(\cuif.ALUOP[3]~4_combout ),
	.datac(\Equal25~0_combout ),
	.datad(Equal0),
	.cin(gnd),
	.combout(\cuif.ALUOP[3]~7_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[3]~7 .lut_mask = 16'h0008;
defparam \cuif.ALUOP[3]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N4
cycloneive_lcell_comb \cuif.ALUOP[3]~5 (
// Equation(s):
// \cuif.ALUOP[3]~5_combout  = (cuifRegWEN & (\cuif.ALUOP[3]~4_combout  & (\Equal25~0_combout  & !Equal0)))

	.dataa(cuifRegWEN),
	.datab(\cuif.ALUOP[3]~4_combout ),
	.datac(\Equal25~0_combout ),
	.datad(Equal0),
	.cin(gnd),
	.combout(\cuif.ALUOP[3]~5_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[3]~5 .lut_mask = 16'h0080;
defparam \cuif.ALUOP[3]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N18
cycloneive_lcell_comb \cuif.ALUOP[3]~6 (
// Equation(s):
// \cuif.ALUOP[3]~6_combout  = (dcifimemload_5 & (dcifimemload_1 & \always0~0_combout ))

	.dataa(gnd),
	.datab(dcifimemload_5),
	.datac(dcifimemload_1),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\cuif.ALUOP[3]~6_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[3]~6 .lut_mask = 16'hC000;
defparam \cuif.ALUOP[3]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N20
cycloneive_lcell_comb \cuif.ALUOP[2]~9 (
// Equation(s):
// \cuif.ALUOP[2]~9_combout  = (dcifimemload_2 & (!dcifimemload_3 & (!dcifimemload_4 & dcifimemload_5)))

	.dataa(dcifimemload_2),
	.datab(dcifimemload_3),
	.datac(dcifimemload_4),
	.datad(dcifimemload_5),
	.cin(gnd),
	.combout(\cuif.ALUOP[2]~9_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[2]~9 .lut_mask = 16'h0200;
defparam \cuif.ALUOP[2]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N26
cycloneive_lcell_comb \cuif.ALUOP[2]~10 (
// Equation(s):
// \cuif.ALUOP[2]~10_combout  = (Equal0 & (\cuif.ALUOP[2]~9_combout )) # (!Equal0 & (((cuifRegWEN & \Equal8~0_combout ))))

	.dataa(Equal0),
	.datab(\cuif.ALUOP[2]~9_combout ),
	.datac(cuifRegWEN),
	.datad(\Equal8~0_combout ),
	.cin(gnd),
	.combout(\cuif.ALUOP[2]~10_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[2]~10 .lut_mask = 16'hD888;
defparam \cuif.ALUOP[2]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N6
cycloneive_lcell_comb \cuif.ALUOP[1]~12 (
// Equation(s):
// \cuif.ALUOP[1]~12_combout  = (dcifimemload_2 & (!dcifimemload_4 & !dcifimemload_3))

	.dataa(dcifimemload_2),
	.datab(gnd),
	.datac(dcifimemload_4),
	.datad(dcifimemload_3),
	.cin(gnd),
	.combout(\cuif.ALUOP[1]~12_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[1]~12 .lut_mask = 16'h000A;
defparam \cuif.ALUOP[1]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N24
cycloneive_lcell_comb \cuif.ALUOP[1]~13 (
// Equation(s):
// \cuif.ALUOP[1]~13_combout  = ((dcifimemload_5 & ((dcifimemload_1))) # (!dcifimemload_5 & (dcifimemload_0))) # (!\cuif.ALUOP[1]~12_combout )

	.dataa(dcifimemload_0),
	.datab(dcifimemload_1),
	.datac(dcifimemload_5),
	.datad(\cuif.ALUOP[1]~12_combout ),
	.cin(gnd),
	.combout(\cuif.ALUOP[1]~13_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[1]~13 .lut_mask = 16'hCAFF;
defparam \cuif.ALUOP[1]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N26
cycloneive_lcell_comb \cuif.ALUOP[1]~14 (
// Equation(s):
// \cuif.ALUOP[1]~14_combout  = (\cuif.ALUOP[1]~3_combout  & ((dcifimemload_28) # ((!dcifimemload_26 & \cuif.ALUOP[1]~13_combout ))))

	.dataa(dcifimemload_26),
	.datab(dcifimemload_28),
	.datac(\cuif.ALUOP[1]~3_combout ),
	.datad(\cuif.ALUOP[1]~13_combout ),
	.cin(gnd),
	.combout(\cuif.ALUOP[1]~14_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[1]~14 .lut_mask = 16'hD0C0;
defparam \cuif.ALUOP[1]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N18
cycloneive_lcell_comb \Equal11~2 (
// Equation(s):
// \Equal11~2_combout  = (Equal3 & ((ccifiwait_0 & (ramiframload_31)) # (!ccifiwait_0 & ((instr_31)))))

	.dataa(ccifiwait_0),
	.datab(Equal3),
	.datac(ramiframload_31),
	.datad(instr_31),
	.cin(gnd),
	.combout(\Equal11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal11~2 .lut_mask = 16'hC480;
defparam \Equal11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N28
cycloneive_lcell_comb \cuif.ALUOP[1]~15 (
// Equation(s):
// \cuif.ALUOP[1]~15_combout  = (dcifimemload_29 & (((!dcifimemload_26 & dcifimemload_27)) # (!dcifimemload_28)))

	.dataa(dcifimemload_26),
	.datab(dcifimemload_29),
	.datac(dcifimemload_27),
	.datad(dcifimemload_28),
	.cin(gnd),
	.combout(\cuif.ALUOP[1]~15_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[1]~15 .lut_mask = 16'h40CC;
defparam \cuif.ALUOP[1]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N10
cycloneive_lcell_comb \cuif.ALUOP[0]~21 (
// Equation(s):
// \cuif.ALUOP[0]~21_combout  = (dcifimemload_2 & (!dcifimemload_3 & (dcifimemload_0 $ (dcifimemload_1)))) # (!dcifimemload_2 & (dcifimemload_0 & (dcifimemload_1 & dcifimemload_3)))

	.dataa(dcifimemload_0),
	.datab(dcifimemload_1),
	.datac(dcifimemload_2),
	.datad(dcifimemload_3),
	.cin(gnd),
	.combout(\cuif.ALUOP[0]~21_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[0]~21 .lut_mask = 16'h0860;
defparam \cuif.ALUOP[0]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N22
cycloneive_lcell_comb \cuif.ALUOP[0]~22 (
// Equation(s):
// \cuif.ALUOP[0]~22_combout  = (dcifimemload_3 & (dcifimemload_1 & (dcifimemload_5 & \cuif.ALUOP[0]~21_combout ))) # (!dcifimemload_3 & ((dcifimemload_1 & (dcifimemload_5 $ (\cuif.ALUOP[0]~21_combout ))) # (!dcifimemload_1 & (dcifimemload_5 & 
// \cuif.ALUOP[0]~21_combout ))))

	.dataa(dcifimemload_3),
	.datab(dcifimemload_1),
	.datac(dcifimemload_5),
	.datad(\cuif.ALUOP[0]~21_combout ),
	.cin(gnd),
	.combout(\cuif.ALUOP[0]~22_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[0]~22 .lut_mask = 16'h9440;
defparam \cuif.ALUOP[0]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N4
cycloneive_lcell_comb \cuif.ALUOP[0]~18 (
// Equation(s):
// \cuif.ALUOP[0]~18_combout  = (!dcifimemload_4 & (\cuif.ALUOP[0]~22_combout  & Equal0))

	.dataa(dcifimemload_4),
	.datab(gnd),
	.datac(\cuif.ALUOP[0]~22_combout ),
	.datad(Equal0),
	.cin(gnd),
	.combout(\cuif.ALUOP[0]~18_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[0]~18 .lut_mask = 16'h5000;
defparam \cuif.ALUOP[0]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N24
cycloneive_lcell_comb \Equal7~1 (
// Equation(s):
// \Equal7~1_combout  = (Equal7 & (dcifimemload_26 & !dcifimemload_27))

	.dataa(Equal7),
	.datab(gnd),
	.datac(dcifimemload_26),
	.datad(dcifimemload_27),
	.cin(gnd),
	.combout(\Equal7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal7~1 .lut_mask = 16'h00A0;
defparam \Equal7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N18
cycloneive_lcell_comb \cuif.ALUOP[0]~17 (
// Equation(s):
// \cuif.ALUOP[0]~17_combout  = (!\Equal25~0_combout  & (!Equal0 & (\Equal7~1_combout  & \cuif.ALUOP[3]~4_combout )))

	.dataa(\Equal25~0_combout ),
	.datab(Equal0),
	.datac(\Equal7~1_combout ),
	.datad(\cuif.ALUOP[3]~4_combout ),
	.cin(gnd),
	.combout(\cuif.ALUOP[0]~17_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.ALUOP[0]~17 .lut_mask = 16'h1000;
defparam \cuif.ALUOP[0]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N24
cycloneive_lcell_comb \Equal4~0 (
// Equation(s):
// \Equal4~0_combout  = (dcifimemload_28 & (\Equal0~1_combout  & \cuif.ALUOP[1]~3_combout ))

	.dataa(dcifimemload_28),
	.datab(\Equal0~1_combout ),
	.datac(gnd),
	.datad(\cuif.ALUOP[1]~3_combout ),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal4~0 .lut_mask = 16'h8800;
defparam \Equal4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N28
cycloneive_lcell_comb \cuif.PCSrc[0]~0 (
// Equation(s):
// \cuif.PCSrc[0]~0_combout  = (\Equal4~0_combout  & (!Equal31 & !Equal2))

	.dataa(\Equal4~0_combout ),
	.datab(Equal31),
	.datac(gnd),
	.datad(Equal2),
	.cin(gnd),
	.combout(\cuif.PCSrc[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.PCSrc[0]~0 .lut_mask = 16'h0022;
defparam \cuif.PCSrc[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N6
cycloneive_lcell_comb \Equal10~0 (
// Equation(s):
// \Equal10~0_combout  = (dcifimemload_27 & (dcifimemload_26 & Equal7))

	.dataa(gnd),
	.datab(dcifimemload_27),
	.datac(dcifimemload_26),
	.datad(Equal7),
	.cin(gnd),
	.combout(\Equal10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~0 .lut_mask = 16'hC000;
defparam \Equal10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N28
cycloneive_lcell_comb \cuif.RegWEN~1 (
// Equation(s):
// \cuif.RegWEN~1_combout  = (!always0 & (((!dcifimemload_29 & dcifdhit)) # (!\Equal11~2_combout )))

	.dataa(\Equal11~2_combout ),
	.datab(dcifimemload_29),
	.datac(dcifdhit),
	.datad(always0),
	.cin(gnd),
	.combout(\cuif.RegWEN~1_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.RegWEN~1 .lut_mask = 16'h0075;
defparam \cuif.RegWEN~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module program_counter_unit (
	PC_29,
	PC_28,
	PC_31,
	PC_30,
	PC_1,
	PC_0,
	PC_3,
	PC_2,
	PC_5,
	PC_4,
	PC_7,
	PC_6,
	PC_9,
	PC_8,
	PC_11,
	PC_10,
	PC_13,
	PC_12,
	PC_15,
	PC_14,
	PC_17,
	PC_16,
	PC_19,
	PC_18,
	PC_21,
	PC_20,
	PC_23,
	PC_22,
	PC_25,
	PC_24,
	PC_27,
	PC_26,
	\pcuif.ihit ,
	dcifimemload_19,
	dcifimemload_18,
	dcifimemload_16,
	dcifimemload_17,
	dcifimemload_20,
	dcifimemload_24,
	dcifimemload_23,
	dcifimemload_21,
	dcifimemload_22,
	Mux30,
	Mux301,
	dcifimemload_25,
	dcifimemload_3,
	dcifimemload_4,
	dcifimemload_2,
	dcifimemload_5,
	dcifimemload_0,
	dcifimemload_1,
	always0,
	Mux0,
	dcifimemload_15,
	Mux1,
	Mux2,
	Mux3,
	Mux4,
	Mux5,
	Mux6,
	Mux7,
	Mux8,
	Mux9,
	Mux10,
	Mux11,
	Mux12,
	Mux13,
	Mux14,
	Mux15,
	Mux16,
	Mux17,
	dcifimemload_14,
	Mux18,
	dcifimemload_13,
	Mux19,
	dcifimemload_12,
	Mux20,
	dcifimemload_11,
	Mux21,
	dcifimemload_10,
	Mux22,
	dcifimemload_9,
	Mux23,
	dcifimemload_8,
	Mux24,
	dcifimemload_7,
	Mux25,
	dcifimemload_6,
	Mux26,
	Mux27,
	Mux28,
	Mux29,
	Mux31,
	Mux311,
	Equal2,
	Equal3,
	cuifPCSrc_0,
	cuifPCSrc_1,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
output 	PC_29;
output 	PC_28;
output 	PC_31;
output 	PC_30;
output 	PC_1;
output 	PC_0;
output 	PC_3;
output 	PC_2;
output 	PC_5;
output 	PC_4;
output 	PC_7;
output 	PC_6;
output 	PC_9;
output 	PC_8;
output 	PC_11;
output 	PC_10;
output 	PC_13;
output 	PC_12;
output 	PC_15;
output 	PC_14;
output 	PC_17;
output 	PC_16;
output 	PC_19;
output 	PC_18;
output 	PC_21;
output 	PC_20;
output 	PC_23;
output 	PC_22;
output 	PC_25;
output 	PC_24;
output 	PC_27;
output 	PC_26;
input 	\pcuif.ihit ;
input 	dcifimemload_19;
input 	dcifimemload_18;
input 	dcifimemload_16;
input 	dcifimemload_17;
input 	dcifimemload_20;
input 	dcifimemload_24;
input 	dcifimemload_23;
input 	dcifimemload_21;
input 	dcifimemload_22;
input 	Mux30;
input 	Mux301;
input 	dcifimemload_25;
input 	dcifimemload_3;
input 	dcifimemload_4;
input 	dcifimemload_2;
input 	dcifimemload_5;
input 	dcifimemload_0;
input 	dcifimemload_1;
input 	always0;
input 	Mux0;
input 	dcifimemload_15;
input 	Mux1;
input 	Mux2;
input 	Mux3;
input 	Mux4;
input 	Mux5;
input 	Mux6;
input 	Mux7;
input 	Mux8;
input 	Mux9;
input 	Mux10;
input 	Mux11;
input 	Mux12;
input 	Mux13;
input 	Mux14;
input 	Mux15;
input 	Mux16;
input 	Mux17;
input 	dcifimemload_14;
input 	Mux18;
input 	dcifimemload_13;
input 	Mux19;
input 	dcifimemload_12;
input 	Mux20;
input 	dcifimemload_11;
input 	Mux21;
input 	dcifimemload_10;
input 	Mux22;
input 	dcifimemload_9;
input 	Mux23;
input 	dcifimemload_8;
input 	Mux24;
input 	dcifimemload_7;
input 	Mux25;
input 	dcifimemload_6;
input 	Mux26;
input 	Mux27;
input 	Mux28;
input 	Mux29;
input 	Mux31;
input 	Mux311;
input 	Equal2;
input 	Equal3;
input 	cuifPCSrc_0;
input 	cuifPCSrc_1;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~2_combout ;
wire \npc[4]~4_combout ;
wire \npc[5]~6_combout ;
wire \Add1~30_combout ;
wire \npc[21]~38_combout ;
wire \npc[24]~44_combout ;
wire \npc[2]~1 ;
wire \npc[3]~3 ;
wire \npc[4]~5 ;
wire \npc[5]~7 ;
wire \npc[6]~9 ;
wire \npc[7]~11 ;
wire \npc[8]~13 ;
wire \npc[9]~15 ;
wire \npc[10]~17 ;
wire \npc[11]~19 ;
wire \npc[12]~21 ;
wire \npc[13]~23 ;
wire \npc[14]~25 ;
wire \npc[15]~27 ;
wire \npc[16]~29 ;
wire \npc[17]~31 ;
wire \npc[18]~33 ;
wire \npc[19]~35 ;
wire \npc[20]~37 ;
wire \npc[21]~39 ;
wire \npc[22]~41 ;
wire \npc[23]~43 ;
wire \npc[24]~45 ;
wire \npc[25]~47 ;
wire \npc[26]~49 ;
wire \npc[27]~51 ;
wire \npc[28]~53 ;
wire \npc[29]~54_combout ;
wire \npc[28]~52_combout ;
wire \npc[27]~50_combout ;
wire \npc[26]~48_combout ;
wire \npc[25]~46_combout ;
wire \npc[23]~42_combout ;
wire \npc[18]~32_combout ;
wire \npc[15]~26_combout ;
wire \npc[13]~22_combout ;
wire \npc[11]~18_combout ;
wire \npc[10]~16_combout ;
wire \npc[7]~10_combout ;
wire \npc[6]~8_combout ;
wire \npc[3]~2_combout ;
wire \npc[2]~0_combout ;
wire \Add1~1 ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~7 ;
wire \Add1~9 ;
wire \Add1~11 ;
wire \Add1~13 ;
wire \Add1~15 ;
wire \Add1~17 ;
wire \Add1~19 ;
wire \Add1~21 ;
wire \Add1~23 ;
wire \Add1~25 ;
wire \Add1~27 ;
wire \Add1~29 ;
wire \Add1~31 ;
wire \Add1~33 ;
wire \Add1~35 ;
wire \Add1~37 ;
wire \Add1~39 ;
wire \Add1~41 ;
wire \Add1~43 ;
wire \Add1~45 ;
wire \Add1~47 ;
wire \Add1~49 ;
wire \Add1~51 ;
wire \Add1~53 ;
wire \Add1~54_combout ;
wire \PC[29]~1_combout ;
wire \Add1~52_combout ;
wire \PC[28]~0_combout ;
wire \npc[29]~55 ;
wire \npc[30]~57 ;
wire \npc[31]~58_combout ;
wire \Add1~55 ;
wire \Add1~57 ;
wire \Add1~58_combout ;
wire \PC[31]~3_combout ;
wire \Add1~56_combout ;
wire \PC[30]~2_combout ;
wire \npc[30]~56_combout ;
wire \Mux30~2_combout ;
wire \PC[1]~4_combout ;
wire \Mux31~2_combout ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \Add1~0_combout ;
wire \Mux29~0_combout ;
wire \Mux29~1_combout ;
wire \Add1~6_combout ;
wire \Mux26~0_combout ;
wire \Mux26~1_combout ;
wire \Add1~4_combout ;
wire \Mux27~0_combout ;
wire \Mux27~1_combout ;
wire \Add1~10_combout ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \Add1~8_combout ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \npc[9]~14_combout ;
wire \Add1~14_combout ;
wire \Mux22~0_combout ;
wire \Mux22~1_combout ;
wire \Add1~12_combout ;
wire \npc[8]~12_combout ;
wire \Mux23~0_combout ;
wire \Mux23~1_combout ;
wire \Add1~18_combout ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \Add1~16_combout ;
wire \Mux21~0_combout ;
wire \Mux21~1_combout ;
wire \Add1~22_combout ;
wire \Mux18~0_combout ;
wire \Mux18~1_combout ;
wire \Add1~20_combout ;
wire \npc[12]~20_combout ;
wire \Mux19~0_combout ;
wire \Mux19~1_combout ;
wire \Add1~26_combout ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \Add1~24_combout ;
wire \npc[14]~24_combout ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \npc[17]~30_combout ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \Add1~28_combout ;
wire \npc[16]~28_combout ;
wire \Mux15~0_combout ;
wire \Mux15~1_combout ;
wire \npc[19]~34_combout ;
wire \Add1~34_combout ;
wire \Mux12~0_combout ;
wire \Mux12~1_combout ;
wire \Add1~32_combout ;
wire \Mux13~0_combout ;
wire \Mux13~1_combout ;
wire \Add1~38_combout ;
wire \Mux10~0_combout ;
wire \Mux10~1_combout ;
wire \Add1~36_combout ;
wire \npc[20]~36_combout ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \Add1~42_combout ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \Add1~40_combout ;
wire \npc[22]~40_combout ;
wire \Mux9~0_combout ;
wire \Mux9~1_combout ;
wire \Add1~46_combout ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \Add1~44_combout ;
wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \Add1~50_combout ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;
wire \Add1~48_combout ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;


// Location: LCCOMB_X61_Y30_N4
cycloneive_lcell_comb \Add1~2 (
// Equation(s):
// \Add1~2_combout  = (dcifimemload_1 & ((\npc[3]~2_combout  & (\Add1~1  & VCC)) # (!\npc[3]~2_combout  & (!\Add1~1 )))) # (!dcifimemload_1 & ((\npc[3]~2_combout  & (!\Add1~1 )) # (!\npc[3]~2_combout  & ((\Add1~1 ) # (GND)))))
// \Add1~3  = CARRY((dcifimemload_1 & (!\npc[3]~2_combout  & !\Add1~1 )) # (!dcifimemload_1 & ((!\Add1~1 ) # (!\npc[3]~2_combout ))))

	.dataa(dcifimemload_1),
	.datab(\npc[3]~2_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h9617;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N6
cycloneive_lcell_comb \npc[4]~4 (
// Equation(s):
// \npc[4]~4_combout  = (PC_4 & (\npc[3]~3  $ (GND))) # (!PC_4 & (!\npc[3]~3  & VCC))
// \npc[4]~5  = CARRY((PC_4 & !\npc[3]~3 ))

	.dataa(gnd),
	.datab(PC_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[3]~3 ),
	.combout(\npc[4]~4_combout ),
	.cout(\npc[4]~5 ));
// synopsys translate_off
defparam \npc[4]~4 .lut_mask = 16'hC30C;
defparam \npc[4]~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N8
cycloneive_lcell_comb \npc[5]~6 (
// Equation(s):
// \npc[5]~6_combout  = (PC_5 & (!\npc[4]~5 )) # (!PC_5 & ((\npc[4]~5 ) # (GND)))
// \npc[5]~7  = CARRY((!\npc[4]~5 ) # (!PC_5))

	.dataa(gnd),
	.datab(PC_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[4]~5 ),
	.combout(\npc[5]~6_combout ),
	.cout(\npc[5]~7 ));
// synopsys translate_off
defparam \npc[5]~6 .lut_mask = 16'h3C3F;
defparam \npc[5]~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N0
cycloneive_lcell_comb \Add1~30 (
// Equation(s):
// \Add1~30_combout  = (\npc[17]~30_combout  & ((dcifimemload_15 & (\Add1~29  & VCC)) # (!dcifimemload_15 & (!\Add1~29 )))) # (!\npc[17]~30_combout  & ((dcifimemload_15 & (!\Add1~29 )) # (!dcifimemload_15 & ((\Add1~29 ) # (GND)))))
// \Add1~31  = CARRY((\npc[17]~30_combout  & (!dcifimemload_15 & !\Add1~29 )) # (!\npc[17]~30_combout  & ((!\Add1~29 ) # (!dcifimemload_15))))

	.dataa(\npc[17]~30_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~29 ),
	.combout(\Add1~30_combout ),
	.cout(\Add1~31 ));
// synopsys translate_off
defparam \Add1~30 .lut_mask = 16'h9617;
defparam \Add1~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N8
cycloneive_lcell_comb \npc[21]~38 (
// Equation(s):
// \npc[21]~38_combout  = (PC_21 & (!\npc[20]~37 )) # (!PC_21 & ((\npc[20]~37 ) # (GND)))
// \npc[21]~39  = CARRY((!\npc[20]~37 ) # (!PC_21))

	.dataa(gnd),
	.datab(PC_21),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[20]~37 ),
	.combout(\npc[21]~38_combout ),
	.cout(\npc[21]~39 ));
// synopsys translate_off
defparam \npc[21]~38 .lut_mask = 16'h3C3F;
defparam \npc[21]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N14
cycloneive_lcell_comb \npc[24]~44 (
// Equation(s):
// \npc[24]~44_combout  = (PC_24 & (\npc[23]~43  $ (GND))) # (!PC_24 & (!\npc[23]~43  & VCC))
// \npc[24]~45  = CARRY((PC_24 & !\npc[23]~43 ))

	.dataa(PC_24),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[23]~43 ),
	.combout(\npc[24]~44_combout ),
	.cout(\npc[24]~45 ));
// synopsys translate_off
defparam \npc[24]~44 .lut_mask = 16'hA50A;
defparam \npc[24]~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X57_Y32_N9
dffeas \PC[29] (
	.clk(CLK),
	.d(\PC[29]~1_combout ),
	.asdata(\npc[29]~54_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(cuifPCSrc_0),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_29),
	.prn(vcc));
// synopsys translate_off
defparam \PC[29] .is_wysiwyg = "true";
defparam \PC[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y29_N17
dffeas \PC[28] (
	.clk(CLK),
	.d(\PC[28]~0_combout ),
	.asdata(\npc[28]~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(cuifPCSrc_0),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_28),
	.prn(vcc));
// synopsys translate_off
defparam \PC[28] .is_wysiwyg = "true";
defparam \PC[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N29
dffeas \PC[31] (
	.clk(CLK),
	.d(\PC[31]~3_combout ),
	.asdata(\npc[31]~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(cuifPCSrc_0),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_31),
	.prn(vcc));
// synopsys translate_off
defparam \PC[31] .is_wysiwyg = "true";
defparam \PC[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y29_N31
dffeas \PC[30] (
	.clk(CLK),
	.d(\PC[30]~2_combout ),
	.asdata(\npc[30]~56_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(cuifPCSrc_0),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_30),
	.prn(vcc));
// synopsys translate_off
defparam \PC[30] .is_wysiwyg = "true";
defparam \PC[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N27
dffeas \PC[1] (
	.clk(CLK),
	.d(\Mux30~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC[1]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_1),
	.prn(vcc));
// synopsys translate_off
defparam \PC[1] .is_wysiwyg = "true";
defparam \PC[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N5
dffeas \PC[0] (
	.clk(CLK),
	.d(\Mux31~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\PC[1]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_0),
	.prn(vcc));
// synopsys translate_off
defparam \PC[0] .is_wysiwyg = "true";
defparam \PC[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N1
dffeas \PC[3] (
	.clk(CLK),
	.d(\Mux28~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_3),
	.prn(vcc));
// synopsys translate_off
defparam \PC[3] .is_wysiwyg = "true";
defparam \PC[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N3
dffeas \PC[2] (
	.clk(CLK),
	.d(\Mux29~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_2),
	.prn(vcc));
// synopsys translate_off
defparam \PC[2] .is_wysiwyg = "true";
defparam \PC[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N13
dffeas \PC[5] (
	.clk(CLK),
	.d(\Mux26~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_5),
	.prn(vcc));
// synopsys translate_off
defparam \PC[5] .is_wysiwyg = "true";
defparam \PC[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N3
dffeas \PC[4] (
	.clk(CLK),
	.d(\Mux27~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_4),
	.prn(vcc));
// synopsys translate_off
defparam \PC[4] .is_wysiwyg = "true";
defparam \PC[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N1
dffeas \PC[7] (
	.clk(CLK),
	.d(\Mux24~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_7),
	.prn(vcc));
// synopsys translate_off
defparam \PC[7] .is_wysiwyg = "true";
defparam \PC[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N5
dffeas \PC[6] (
	.clk(CLK),
	.d(\Mux25~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_6),
	.prn(vcc));
// synopsys translate_off
defparam \PC[6] .is_wysiwyg = "true";
defparam \PC[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N31
dffeas \PC[9] (
	.clk(CLK),
	.d(\Mux22~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_9),
	.prn(vcc));
// synopsys translate_off
defparam \PC[9] .is_wysiwyg = "true";
defparam \PC[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N9
dffeas \PC[8] (
	.clk(CLK),
	.d(\Mux23~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_8),
	.prn(vcc));
// synopsys translate_off
defparam \PC[8] .is_wysiwyg = "true";
defparam \PC[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N13
dffeas \PC[11] (
	.clk(CLK),
	.d(\Mux20~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_11),
	.prn(vcc));
// synopsys translate_off
defparam \PC[11] .is_wysiwyg = "true";
defparam \PC[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N31
dffeas \PC[10] (
	.clk(CLK),
	.d(\Mux21~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_10),
	.prn(vcc));
// synopsys translate_off
defparam \PC[10] .is_wysiwyg = "true";
defparam \PC[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N5
dffeas \PC[13] (
	.clk(CLK),
	.d(\Mux18~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_13),
	.prn(vcc));
// synopsys translate_off
defparam \PC[13] .is_wysiwyg = "true";
defparam \PC[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N23
dffeas \PC[12] (
	.clk(CLK),
	.d(\Mux19~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_12),
	.prn(vcc));
// synopsys translate_off
defparam \PC[12] .is_wysiwyg = "true";
defparam \PC[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N21
dffeas \PC[15] (
	.clk(CLK),
	.d(\Mux16~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_15),
	.prn(vcc));
// synopsys translate_off
defparam \PC[15] .is_wysiwyg = "true";
defparam \PC[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N15
dffeas \PC[14] (
	.clk(CLK),
	.d(\Mux17~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_14),
	.prn(vcc));
// synopsys translate_off
defparam \PC[14] .is_wysiwyg = "true";
defparam \PC[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N1
dffeas \PC[17] (
	.clk(CLK),
	.d(\Mux14~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_17),
	.prn(vcc));
// synopsys translate_off
defparam \PC[17] .is_wysiwyg = "true";
defparam \PC[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N1
dffeas \PC[16] (
	.clk(CLK),
	.d(\Mux15~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_16),
	.prn(vcc));
// synopsys translate_off
defparam \PC[16] .is_wysiwyg = "true";
defparam \PC[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N11
dffeas \PC[19] (
	.clk(CLK),
	.d(\Mux12~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_19),
	.prn(vcc));
// synopsys translate_off
defparam \PC[19] .is_wysiwyg = "true";
defparam \PC[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N29
dffeas \PC[18] (
	.clk(CLK),
	.d(\Mux13~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_18),
	.prn(vcc));
// synopsys translate_off
defparam \PC[18] .is_wysiwyg = "true";
defparam \PC[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N21
dffeas \PC[21] (
	.clk(CLK),
	.d(\Mux10~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_21),
	.prn(vcc));
// synopsys translate_off
defparam \PC[21] .is_wysiwyg = "true";
defparam \PC[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N3
dffeas \PC[20] (
	.clk(CLK),
	.d(\Mux11~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_20),
	.prn(vcc));
// synopsys translate_off
defparam \PC[20] .is_wysiwyg = "true";
defparam \PC[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N5
dffeas \PC[23] (
	.clk(CLK),
	.d(\Mux8~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_23),
	.prn(vcc));
// synopsys translate_off
defparam \PC[23] .is_wysiwyg = "true";
defparam \PC[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N17
dffeas \PC[22] (
	.clk(CLK),
	.d(\Mux9~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_22),
	.prn(vcc));
// synopsys translate_off
defparam \PC[22] .is_wysiwyg = "true";
defparam \PC[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N9
dffeas \PC[25] (
	.clk(CLK),
	.d(\Mux6~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_25),
	.prn(vcc));
// synopsys translate_off
defparam \PC[25] .is_wysiwyg = "true";
defparam \PC[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N31
dffeas \PC[24] (
	.clk(CLK),
	.d(\Mux7~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_24),
	.prn(vcc));
// synopsys translate_off
defparam \PC[24] .is_wysiwyg = "true";
defparam \PC[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N13
dffeas \PC[27] (
	.clk(CLK),
	.d(\Mux4~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_27),
	.prn(vcc));
// synopsys translate_off
defparam \PC[27] .is_wysiwyg = "true";
defparam \PC[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N25
dffeas \PC[26] (
	.clk(CLK),
	.d(\Mux5~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcuif.ihit ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PC_26),
	.prn(vcc));
// synopsys translate_off
defparam \PC[26] .is_wysiwyg = "true";
defparam \PC[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N2
cycloneive_lcell_comb \npc[2]~0 (
// Equation(s):
// \npc[2]~0_combout  = PC_2 $ (VCC)
// \npc[2]~1  = CARRY(PC_2)

	.dataa(gnd),
	.datab(PC_2),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\npc[2]~0_combout ),
	.cout(\npc[2]~1 ));
// synopsys translate_off
defparam \npc[2]~0 .lut_mask = 16'h33CC;
defparam \npc[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N4
cycloneive_lcell_comb \npc[3]~2 (
// Equation(s):
// \npc[3]~2_combout  = (PC_3 & (!\npc[2]~1 )) # (!PC_3 & ((\npc[2]~1 ) # (GND)))
// \npc[3]~3  = CARRY((!\npc[2]~1 ) # (!PC_3))

	.dataa(PC_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[2]~1 ),
	.combout(\npc[3]~2_combout ),
	.cout(\npc[3]~3 ));
// synopsys translate_off
defparam \npc[3]~2 .lut_mask = 16'h5A5F;
defparam \npc[3]~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N10
cycloneive_lcell_comb \npc[6]~8 (
// Equation(s):
// \npc[6]~8_combout  = (PC_6 & (\npc[5]~7  $ (GND))) # (!PC_6 & (!\npc[5]~7  & VCC))
// \npc[6]~9  = CARRY((PC_6 & !\npc[5]~7 ))

	.dataa(gnd),
	.datab(PC_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[5]~7 ),
	.combout(\npc[6]~8_combout ),
	.cout(\npc[6]~9 ));
// synopsys translate_off
defparam \npc[6]~8 .lut_mask = 16'hC30C;
defparam \npc[6]~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N12
cycloneive_lcell_comb \npc[7]~10 (
// Equation(s):
// \npc[7]~10_combout  = (PC_7 & (!\npc[6]~9 )) # (!PC_7 & ((\npc[6]~9 ) # (GND)))
// \npc[7]~11  = CARRY((!\npc[6]~9 ) # (!PC_7))

	.dataa(PC_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[6]~9 ),
	.combout(\npc[7]~10_combout ),
	.cout(\npc[7]~11 ));
// synopsys translate_off
defparam \npc[7]~10 .lut_mask = 16'h5A5F;
defparam \npc[7]~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N14
cycloneive_lcell_comb \npc[8]~12 (
// Equation(s):
// \npc[8]~12_combout  = (PC_8 & (\npc[7]~11  $ (GND))) # (!PC_8 & (!\npc[7]~11  & VCC))
// \npc[8]~13  = CARRY((PC_8 & !\npc[7]~11 ))

	.dataa(PC_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[7]~11 ),
	.combout(\npc[8]~12_combout ),
	.cout(\npc[8]~13 ));
// synopsys translate_off
defparam \npc[8]~12 .lut_mask = 16'hA50A;
defparam \npc[8]~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N16
cycloneive_lcell_comb \npc[9]~14 (
// Equation(s):
// \npc[9]~14_combout  = (PC_9 & (!\npc[8]~13 )) # (!PC_9 & ((\npc[8]~13 ) # (GND)))
// \npc[9]~15  = CARRY((!\npc[8]~13 ) # (!PC_9))

	.dataa(gnd),
	.datab(PC_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[8]~13 ),
	.combout(\npc[9]~14_combout ),
	.cout(\npc[9]~15 ));
// synopsys translate_off
defparam \npc[9]~14 .lut_mask = 16'h3C3F;
defparam \npc[9]~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N18
cycloneive_lcell_comb \npc[10]~16 (
// Equation(s):
// \npc[10]~16_combout  = (PC_10 & (\npc[9]~15  $ (GND))) # (!PC_10 & (!\npc[9]~15  & VCC))
// \npc[10]~17  = CARRY((PC_10 & !\npc[9]~15 ))

	.dataa(gnd),
	.datab(PC_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[9]~15 ),
	.combout(\npc[10]~16_combout ),
	.cout(\npc[10]~17 ));
// synopsys translate_off
defparam \npc[10]~16 .lut_mask = 16'hC30C;
defparam \npc[10]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N20
cycloneive_lcell_comb \npc[11]~18 (
// Equation(s):
// \npc[11]~18_combout  = (PC_11 & (!\npc[10]~17 )) # (!PC_11 & ((\npc[10]~17 ) # (GND)))
// \npc[11]~19  = CARRY((!\npc[10]~17 ) # (!PC_11))

	.dataa(PC_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[10]~17 ),
	.combout(\npc[11]~18_combout ),
	.cout(\npc[11]~19 ));
// synopsys translate_off
defparam \npc[11]~18 .lut_mask = 16'h5A5F;
defparam \npc[11]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N22
cycloneive_lcell_comb \npc[12]~20 (
// Equation(s):
// \npc[12]~20_combout  = (PC_12 & (\npc[11]~19  $ (GND))) # (!PC_12 & (!\npc[11]~19  & VCC))
// \npc[12]~21  = CARRY((PC_12 & !\npc[11]~19 ))

	.dataa(gnd),
	.datab(PC_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[11]~19 ),
	.combout(\npc[12]~20_combout ),
	.cout(\npc[12]~21 ));
// synopsys translate_off
defparam \npc[12]~20 .lut_mask = 16'hC30C;
defparam \npc[12]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N24
cycloneive_lcell_comb \npc[13]~22 (
// Equation(s):
// \npc[13]~22_combout  = (PC_13 & (!\npc[12]~21 )) # (!PC_13 & ((\npc[12]~21 ) # (GND)))
// \npc[13]~23  = CARRY((!\npc[12]~21 ) # (!PC_13))

	.dataa(gnd),
	.datab(PC_13),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[12]~21 ),
	.combout(\npc[13]~22_combout ),
	.cout(\npc[13]~23 ));
// synopsys translate_off
defparam \npc[13]~22 .lut_mask = 16'h3C3F;
defparam \npc[13]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N26
cycloneive_lcell_comb \npc[14]~24 (
// Equation(s):
// \npc[14]~24_combout  = (PC_14 & (\npc[13]~23  $ (GND))) # (!PC_14 & (!\npc[13]~23  & VCC))
// \npc[14]~25  = CARRY((PC_14 & !\npc[13]~23 ))

	.dataa(gnd),
	.datab(PC_14),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[13]~23 ),
	.combout(\npc[14]~24_combout ),
	.cout(\npc[14]~25 ));
// synopsys translate_off
defparam \npc[14]~24 .lut_mask = 16'hC30C;
defparam \npc[14]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N28
cycloneive_lcell_comb \npc[15]~26 (
// Equation(s):
// \npc[15]~26_combout  = (PC_15 & (!\npc[14]~25 )) # (!PC_15 & ((\npc[14]~25 ) # (GND)))
// \npc[15]~27  = CARRY((!\npc[14]~25 ) # (!PC_15))

	.dataa(PC_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[14]~25 ),
	.combout(\npc[15]~26_combout ),
	.cout(\npc[15]~27 ));
// synopsys translate_off
defparam \npc[15]~26 .lut_mask = 16'h5A5F;
defparam \npc[15]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N30
cycloneive_lcell_comb \npc[16]~28 (
// Equation(s):
// \npc[16]~28_combout  = (PC_16 & (\npc[15]~27  $ (GND))) # (!PC_16 & (!\npc[15]~27  & VCC))
// \npc[16]~29  = CARRY((PC_16 & !\npc[15]~27 ))

	.dataa(gnd),
	.datab(PC_16),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[15]~27 ),
	.combout(\npc[16]~28_combout ),
	.cout(\npc[16]~29 ));
// synopsys translate_off
defparam \npc[16]~28 .lut_mask = 16'hC30C;
defparam \npc[16]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N0
cycloneive_lcell_comb \npc[17]~30 (
// Equation(s):
// \npc[17]~30_combout  = (PC_17 & (!\npc[16]~29 )) # (!PC_17 & ((\npc[16]~29 ) # (GND)))
// \npc[17]~31  = CARRY((!\npc[16]~29 ) # (!PC_17))

	.dataa(PC_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[16]~29 ),
	.combout(\npc[17]~30_combout ),
	.cout(\npc[17]~31 ));
// synopsys translate_off
defparam \npc[17]~30 .lut_mask = 16'h5A5F;
defparam \npc[17]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N2
cycloneive_lcell_comb \npc[18]~32 (
// Equation(s):
// \npc[18]~32_combout  = (PC_18 & (\npc[17]~31  $ (GND))) # (!PC_18 & (!\npc[17]~31  & VCC))
// \npc[18]~33  = CARRY((PC_18 & !\npc[17]~31 ))

	.dataa(PC_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[17]~31 ),
	.combout(\npc[18]~32_combout ),
	.cout(\npc[18]~33 ));
// synopsys translate_off
defparam \npc[18]~32 .lut_mask = 16'hA50A;
defparam \npc[18]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N4
cycloneive_lcell_comb \npc[19]~34 (
// Equation(s):
// \npc[19]~34_combout  = (PC_19 & (!\npc[18]~33 )) # (!PC_19 & ((\npc[18]~33 ) # (GND)))
// \npc[19]~35  = CARRY((!\npc[18]~33 ) # (!PC_19))

	.dataa(gnd),
	.datab(PC_19),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[18]~33 ),
	.combout(\npc[19]~34_combout ),
	.cout(\npc[19]~35 ));
// synopsys translate_off
defparam \npc[19]~34 .lut_mask = 16'h3C3F;
defparam \npc[19]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N6
cycloneive_lcell_comb \npc[20]~36 (
// Equation(s):
// \npc[20]~36_combout  = (PC_20 & (\npc[19]~35  $ (GND))) # (!PC_20 & (!\npc[19]~35  & VCC))
// \npc[20]~37  = CARRY((PC_20 & !\npc[19]~35 ))

	.dataa(PC_20),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[19]~35 ),
	.combout(\npc[20]~36_combout ),
	.cout(\npc[20]~37 ));
// synopsys translate_off
defparam \npc[20]~36 .lut_mask = 16'hA50A;
defparam \npc[20]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N10
cycloneive_lcell_comb \npc[22]~40 (
// Equation(s):
// \npc[22]~40_combout  = (PC_22 & (\npc[21]~39  $ (GND))) # (!PC_22 & (!\npc[21]~39  & VCC))
// \npc[22]~41  = CARRY((PC_22 & !\npc[21]~39 ))

	.dataa(gnd),
	.datab(PC_22),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[21]~39 ),
	.combout(\npc[22]~40_combout ),
	.cout(\npc[22]~41 ));
// synopsys translate_off
defparam \npc[22]~40 .lut_mask = 16'hC30C;
defparam \npc[22]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N12
cycloneive_lcell_comb \npc[23]~42 (
// Equation(s):
// \npc[23]~42_combout  = (PC_23 & (!\npc[22]~41 )) # (!PC_23 & ((\npc[22]~41 ) # (GND)))
// \npc[23]~43  = CARRY((!\npc[22]~41 ) # (!PC_23))

	.dataa(gnd),
	.datab(PC_23),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[22]~41 ),
	.combout(\npc[23]~42_combout ),
	.cout(\npc[23]~43 ));
// synopsys translate_off
defparam \npc[23]~42 .lut_mask = 16'h3C3F;
defparam \npc[23]~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N16
cycloneive_lcell_comb \npc[25]~46 (
// Equation(s):
// \npc[25]~46_combout  = (PC_25 & (!\npc[24]~45 )) # (!PC_25 & ((\npc[24]~45 ) # (GND)))
// \npc[25]~47  = CARRY((!\npc[24]~45 ) # (!PC_25))

	.dataa(gnd),
	.datab(PC_25),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[24]~45 ),
	.combout(\npc[25]~46_combout ),
	.cout(\npc[25]~47 ));
// synopsys translate_off
defparam \npc[25]~46 .lut_mask = 16'h3C3F;
defparam \npc[25]~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N18
cycloneive_lcell_comb \npc[26]~48 (
// Equation(s):
// \npc[26]~48_combout  = (PC_26 & (\npc[25]~47  $ (GND))) # (!PC_26 & (!\npc[25]~47  & VCC))
// \npc[26]~49  = CARRY((PC_26 & !\npc[25]~47 ))

	.dataa(gnd),
	.datab(PC_26),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[25]~47 ),
	.combout(\npc[26]~48_combout ),
	.cout(\npc[26]~49 ));
// synopsys translate_off
defparam \npc[26]~48 .lut_mask = 16'hC30C;
defparam \npc[26]~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N20
cycloneive_lcell_comb \npc[27]~50 (
// Equation(s):
// \npc[27]~50_combout  = (PC_27 & (!\npc[26]~49 )) # (!PC_27 & ((\npc[26]~49 ) # (GND)))
// \npc[27]~51  = CARRY((!\npc[26]~49 ) # (!PC_27))

	.dataa(PC_27),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[26]~49 ),
	.combout(\npc[27]~50_combout ),
	.cout(\npc[27]~51 ));
// synopsys translate_off
defparam \npc[27]~50 .lut_mask = 16'h5A5F;
defparam \npc[27]~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N22
cycloneive_lcell_comb \npc[28]~52 (
// Equation(s):
// \npc[28]~52_combout  = (PC_28 & (\npc[27]~51  $ (GND))) # (!PC_28 & (!\npc[27]~51  & VCC))
// \npc[28]~53  = CARRY((PC_28 & !\npc[27]~51 ))

	.dataa(PC_28),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[27]~51 ),
	.combout(\npc[28]~52_combout ),
	.cout(\npc[28]~53 ));
// synopsys translate_off
defparam \npc[28]~52 .lut_mask = 16'hA50A;
defparam \npc[28]~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N24
cycloneive_lcell_comb \npc[29]~54 (
// Equation(s):
// \npc[29]~54_combout  = (PC_29 & (!\npc[28]~53 )) # (!PC_29 & ((\npc[28]~53 ) # (GND)))
// \npc[29]~55  = CARRY((!\npc[28]~53 ) # (!PC_29))

	.dataa(PC_29),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[28]~53 ),
	.combout(\npc[29]~54_combout ),
	.cout(\npc[29]~55 ));
// synopsys translate_off
defparam \npc[29]~54 .lut_mask = 16'h5A5F;
defparam \npc[29]~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N2
cycloneive_lcell_comb \Add1~0 (
// Equation(s):
// \Add1~0_combout  = (dcifimemload_0 & (\npc[2]~0_combout  $ (VCC))) # (!dcifimemload_0 & (\npc[2]~0_combout  & VCC))
// \Add1~1  = CARRY((dcifimemload_0 & \npc[2]~0_combout ))

	.dataa(dcifimemload_0),
	.datab(\npc[2]~0_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h6688;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N6
cycloneive_lcell_comb \Add1~4 (
// Equation(s):
// \Add1~4_combout  = ((\npc[4]~4_combout  $ (dcifimemload_2 $ (!\Add1~3 )))) # (GND)
// \Add1~5  = CARRY((\npc[4]~4_combout  & ((dcifimemload_2) # (!\Add1~3 ))) # (!\npc[4]~4_combout  & (dcifimemload_2 & !\Add1~3 )))

	.dataa(\npc[4]~4_combout ),
	.datab(dcifimemload_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'h698E;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N8
cycloneive_lcell_comb \Add1~6 (
// Equation(s):
// \Add1~6_combout  = (\npc[5]~6_combout  & ((dcifimemload_3 & (\Add1~5  & VCC)) # (!dcifimemload_3 & (!\Add1~5 )))) # (!\npc[5]~6_combout  & ((dcifimemload_3 & (!\Add1~5 )) # (!dcifimemload_3 & ((\Add1~5 ) # (GND)))))
// \Add1~7  = CARRY((\npc[5]~6_combout  & (!dcifimemload_3 & !\Add1~5 )) # (!\npc[5]~6_combout  & ((!\Add1~5 ) # (!dcifimemload_3))))

	.dataa(\npc[5]~6_combout ),
	.datab(dcifimemload_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h9617;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N10
cycloneive_lcell_comb \Add1~8 (
// Equation(s):
// \Add1~8_combout  = ((dcifimemload_4 $ (\npc[6]~8_combout  $ (!\Add1~7 )))) # (GND)
// \Add1~9  = CARRY((dcifimemload_4 & ((\npc[6]~8_combout ) # (!\Add1~7 ))) # (!dcifimemload_4 & (\npc[6]~8_combout  & !\Add1~7 )))

	.dataa(dcifimemload_4),
	.datab(\npc[6]~8_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'h698E;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N12
cycloneive_lcell_comb \Add1~10 (
// Equation(s):
// \Add1~10_combout  = (dcifimemload_5 & ((\npc[7]~10_combout  & (\Add1~9  & VCC)) # (!\npc[7]~10_combout  & (!\Add1~9 )))) # (!dcifimemload_5 & ((\npc[7]~10_combout  & (!\Add1~9 )) # (!\npc[7]~10_combout  & ((\Add1~9 ) # (GND)))))
// \Add1~11  = CARRY((dcifimemload_5 & (!\npc[7]~10_combout  & !\Add1~9 )) # (!dcifimemload_5 & ((!\Add1~9 ) # (!\npc[7]~10_combout ))))

	.dataa(dcifimemload_5),
	.datab(\npc[7]~10_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h9617;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N14
cycloneive_lcell_comb \Add1~12 (
// Equation(s):
// \Add1~12_combout  = ((\npc[8]~12_combout  $ (dcifimemload_6 $ (!\Add1~11 )))) # (GND)
// \Add1~13  = CARRY((\npc[8]~12_combout  & ((dcifimemload_6) # (!\Add1~11 ))) # (!\npc[8]~12_combout  & (dcifimemload_6 & !\Add1~11 )))

	.dataa(\npc[8]~12_combout ),
	.datab(dcifimemload_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
// synopsys translate_off
defparam \Add1~12 .lut_mask = 16'h698E;
defparam \Add1~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N16
cycloneive_lcell_comb \Add1~14 (
// Equation(s):
// \Add1~14_combout  = (\npc[9]~14_combout  & ((dcifimemload_7 & (\Add1~13  & VCC)) # (!dcifimemload_7 & (!\Add1~13 )))) # (!\npc[9]~14_combout  & ((dcifimemload_7 & (!\Add1~13 )) # (!dcifimemload_7 & ((\Add1~13 ) # (GND)))))
// \Add1~15  = CARRY((\npc[9]~14_combout  & (!dcifimemload_7 & !\Add1~13 )) # (!\npc[9]~14_combout  & ((!\Add1~13 ) # (!dcifimemload_7))))

	.dataa(\npc[9]~14_combout ),
	.datab(dcifimemload_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
// synopsys translate_off
defparam \Add1~14 .lut_mask = 16'h9617;
defparam \Add1~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N18
cycloneive_lcell_comb \Add1~16 (
// Equation(s):
// \Add1~16_combout  = ((dcifimemload_8 $ (\npc[10]~16_combout  $ (!\Add1~15 )))) # (GND)
// \Add1~17  = CARRY((dcifimemload_8 & ((\npc[10]~16_combout ) # (!\Add1~15 ))) # (!dcifimemload_8 & (\npc[10]~16_combout  & !\Add1~15 )))

	.dataa(dcifimemload_8),
	.datab(\npc[10]~16_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout(\Add1~17 ));
// synopsys translate_off
defparam \Add1~16 .lut_mask = 16'h698E;
defparam \Add1~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N20
cycloneive_lcell_comb \Add1~18 (
// Equation(s):
// \Add1~18_combout  = (dcifimemload_9 & ((\npc[11]~18_combout  & (\Add1~17  & VCC)) # (!\npc[11]~18_combout  & (!\Add1~17 )))) # (!dcifimemload_9 & ((\npc[11]~18_combout  & (!\Add1~17 )) # (!\npc[11]~18_combout  & ((\Add1~17 ) # (GND)))))
// \Add1~19  = CARRY((dcifimemload_9 & (!\npc[11]~18_combout  & !\Add1~17 )) # (!dcifimemload_9 & ((!\Add1~17 ) # (!\npc[11]~18_combout ))))

	.dataa(dcifimemload_9),
	.datab(\npc[11]~18_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~17 ),
	.combout(\Add1~18_combout ),
	.cout(\Add1~19 ));
// synopsys translate_off
defparam \Add1~18 .lut_mask = 16'h9617;
defparam \Add1~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N22
cycloneive_lcell_comb \Add1~20 (
// Equation(s):
// \Add1~20_combout  = ((\npc[12]~20_combout  $ (dcifimemload_10 $ (!\Add1~19 )))) # (GND)
// \Add1~21  = CARRY((\npc[12]~20_combout  & ((dcifimemload_10) # (!\Add1~19 ))) # (!\npc[12]~20_combout  & (dcifimemload_10 & !\Add1~19 )))

	.dataa(\npc[12]~20_combout ),
	.datab(dcifimemload_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~19 ),
	.combout(\Add1~20_combout ),
	.cout(\Add1~21 ));
// synopsys translate_off
defparam \Add1~20 .lut_mask = 16'h698E;
defparam \Add1~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N24
cycloneive_lcell_comb \Add1~22 (
// Equation(s):
// \Add1~22_combout  = (dcifimemload_11 & ((\npc[13]~22_combout  & (\Add1~21  & VCC)) # (!\npc[13]~22_combout  & (!\Add1~21 )))) # (!dcifimemload_11 & ((\npc[13]~22_combout  & (!\Add1~21 )) # (!\npc[13]~22_combout  & ((\Add1~21 ) # (GND)))))
// \Add1~23  = CARRY((dcifimemload_11 & (!\npc[13]~22_combout  & !\Add1~21 )) # (!dcifimemload_11 & ((!\Add1~21 ) # (!\npc[13]~22_combout ))))

	.dataa(dcifimemload_11),
	.datab(\npc[13]~22_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~21 ),
	.combout(\Add1~22_combout ),
	.cout(\Add1~23 ));
// synopsys translate_off
defparam \Add1~22 .lut_mask = 16'h9617;
defparam \Add1~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N26
cycloneive_lcell_comb \Add1~24 (
// Equation(s):
// \Add1~24_combout  = ((\npc[14]~24_combout  $ (dcifimemload_12 $ (!\Add1~23 )))) # (GND)
// \Add1~25  = CARRY((\npc[14]~24_combout  & ((dcifimemload_12) # (!\Add1~23 ))) # (!\npc[14]~24_combout  & (dcifimemload_12 & !\Add1~23 )))

	.dataa(\npc[14]~24_combout ),
	.datab(dcifimemload_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~23 ),
	.combout(\Add1~24_combout ),
	.cout(\Add1~25 ));
// synopsys translate_off
defparam \Add1~24 .lut_mask = 16'h698E;
defparam \Add1~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N28
cycloneive_lcell_comb \Add1~26 (
// Equation(s):
// \Add1~26_combout  = (dcifimemload_13 & ((\npc[15]~26_combout  & (\Add1~25  & VCC)) # (!\npc[15]~26_combout  & (!\Add1~25 )))) # (!dcifimemload_13 & ((\npc[15]~26_combout  & (!\Add1~25 )) # (!\npc[15]~26_combout  & ((\Add1~25 ) # (GND)))))
// \Add1~27  = CARRY((dcifimemload_13 & (!\npc[15]~26_combout  & !\Add1~25 )) # (!dcifimemload_13 & ((!\Add1~25 ) # (!\npc[15]~26_combout ))))

	.dataa(dcifimemload_13),
	.datab(\npc[15]~26_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~25 ),
	.combout(\Add1~26_combout ),
	.cout(\Add1~27 ));
// synopsys translate_off
defparam \Add1~26 .lut_mask = 16'h9617;
defparam \Add1~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N30
cycloneive_lcell_comb \Add1~28 (
// Equation(s):
// \Add1~28_combout  = ((\npc[16]~28_combout  $ (dcifimemload_14 $ (!\Add1~27 )))) # (GND)
// \Add1~29  = CARRY((\npc[16]~28_combout  & ((dcifimemload_14) # (!\Add1~27 ))) # (!\npc[16]~28_combout  & (dcifimemload_14 & !\Add1~27 )))

	.dataa(\npc[16]~28_combout ),
	.datab(dcifimemload_14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~27 ),
	.combout(\Add1~28_combout ),
	.cout(\Add1~29 ));
// synopsys translate_off
defparam \Add1~28 .lut_mask = 16'h698E;
defparam \Add1~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N2
cycloneive_lcell_comb \Add1~32 (
// Equation(s):
// \Add1~32_combout  = ((dcifimemload_15 $ (\npc[18]~32_combout  $ (!\Add1~31 )))) # (GND)
// \Add1~33  = CARRY((dcifimemload_15 & ((\npc[18]~32_combout ) # (!\Add1~31 ))) # (!dcifimemload_15 & (\npc[18]~32_combout  & !\Add1~31 )))

	.dataa(dcifimemload_15),
	.datab(\npc[18]~32_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~31 ),
	.combout(\Add1~32_combout ),
	.cout(\Add1~33 ));
// synopsys translate_off
defparam \Add1~32 .lut_mask = 16'h698E;
defparam \Add1~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N4
cycloneive_lcell_comb \Add1~34 (
// Equation(s):
// \Add1~34_combout  = (\npc[19]~34_combout  & ((dcifimemload_15 & (\Add1~33  & VCC)) # (!dcifimemload_15 & (!\Add1~33 )))) # (!\npc[19]~34_combout  & ((dcifimemload_15 & (!\Add1~33 )) # (!dcifimemload_15 & ((\Add1~33 ) # (GND)))))
// \Add1~35  = CARRY((\npc[19]~34_combout  & (!dcifimemload_15 & !\Add1~33 )) # (!\npc[19]~34_combout  & ((!\Add1~33 ) # (!dcifimemload_15))))

	.dataa(\npc[19]~34_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~33 ),
	.combout(\Add1~34_combout ),
	.cout(\Add1~35 ));
// synopsys translate_off
defparam \Add1~34 .lut_mask = 16'h9617;
defparam \Add1~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N6
cycloneive_lcell_comb \Add1~36 (
// Equation(s):
// \Add1~36_combout  = ((\npc[20]~36_combout  $ (dcifimemload_15 $ (!\Add1~35 )))) # (GND)
// \Add1~37  = CARRY((\npc[20]~36_combout  & ((dcifimemload_15) # (!\Add1~35 ))) # (!\npc[20]~36_combout  & (dcifimemload_15 & !\Add1~35 )))

	.dataa(\npc[20]~36_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~35 ),
	.combout(\Add1~36_combout ),
	.cout(\Add1~37 ));
// synopsys translate_off
defparam \Add1~36 .lut_mask = 16'h698E;
defparam \Add1~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N8
cycloneive_lcell_comb \Add1~38 (
// Equation(s):
// \Add1~38_combout  = (\npc[21]~38_combout  & ((dcifimemload_15 & (\Add1~37  & VCC)) # (!dcifimemload_15 & (!\Add1~37 )))) # (!\npc[21]~38_combout  & ((dcifimemload_15 & (!\Add1~37 )) # (!dcifimemload_15 & ((\Add1~37 ) # (GND)))))
// \Add1~39  = CARRY((\npc[21]~38_combout  & (!dcifimemload_15 & !\Add1~37 )) # (!\npc[21]~38_combout  & ((!\Add1~37 ) # (!dcifimemload_15))))

	.dataa(\npc[21]~38_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~37 ),
	.combout(\Add1~38_combout ),
	.cout(\Add1~39 ));
// synopsys translate_off
defparam \Add1~38 .lut_mask = 16'h9617;
defparam \Add1~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N10
cycloneive_lcell_comb \Add1~40 (
// Equation(s):
// \Add1~40_combout  = ((\npc[22]~40_combout  $ (dcifimemload_15 $ (!\Add1~39 )))) # (GND)
// \Add1~41  = CARRY((\npc[22]~40_combout  & ((dcifimemload_15) # (!\Add1~39 ))) # (!\npc[22]~40_combout  & (dcifimemload_15 & !\Add1~39 )))

	.dataa(\npc[22]~40_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~39 ),
	.combout(\Add1~40_combout ),
	.cout(\Add1~41 ));
// synopsys translate_off
defparam \Add1~40 .lut_mask = 16'h698E;
defparam \Add1~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N12
cycloneive_lcell_comb \Add1~42 (
// Equation(s):
// \Add1~42_combout  = (dcifimemload_15 & ((\npc[23]~42_combout  & (\Add1~41  & VCC)) # (!\npc[23]~42_combout  & (!\Add1~41 )))) # (!dcifimemload_15 & ((\npc[23]~42_combout  & (!\Add1~41 )) # (!\npc[23]~42_combout  & ((\Add1~41 ) # (GND)))))
// \Add1~43  = CARRY((dcifimemload_15 & (!\npc[23]~42_combout  & !\Add1~41 )) # (!dcifimemload_15 & ((!\Add1~41 ) # (!\npc[23]~42_combout ))))

	.dataa(dcifimemload_15),
	.datab(\npc[23]~42_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~41 ),
	.combout(\Add1~42_combout ),
	.cout(\Add1~43 ));
// synopsys translate_off
defparam \Add1~42 .lut_mask = 16'h9617;
defparam \Add1~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N14
cycloneive_lcell_comb \Add1~44 (
// Equation(s):
// \Add1~44_combout  = ((\npc[24]~44_combout  $ (dcifimemload_15 $ (!\Add1~43 )))) # (GND)
// \Add1~45  = CARRY((\npc[24]~44_combout  & ((dcifimemload_15) # (!\Add1~43 ))) # (!\npc[24]~44_combout  & (dcifimemload_15 & !\Add1~43 )))

	.dataa(\npc[24]~44_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~43 ),
	.combout(\Add1~44_combout ),
	.cout(\Add1~45 ));
// synopsys translate_off
defparam \Add1~44 .lut_mask = 16'h698E;
defparam \Add1~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N16
cycloneive_lcell_comb \Add1~46 (
// Equation(s):
// \Add1~46_combout  = (dcifimemload_15 & ((\npc[25]~46_combout  & (\Add1~45  & VCC)) # (!\npc[25]~46_combout  & (!\Add1~45 )))) # (!dcifimemload_15 & ((\npc[25]~46_combout  & (!\Add1~45 )) # (!\npc[25]~46_combout  & ((\Add1~45 ) # (GND)))))
// \Add1~47  = CARRY((dcifimemload_15 & (!\npc[25]~46_combout  & !\Add1~45 )) # (!dcifimemload_15 & ((!\Add1~45 ) # (!\npc[25]~46_combout ))))

	.dataa(dcifimemload_15),
	.datab(\npc[25]~46_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~45 ),
	.combout(\Add1~46_combout ),
	.cout(\Add1~47 ));
// synopsys translate_off
defparam \Add1~46 .lut_mask = 16'h9617;
defparam \Add1~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N18
cycloneive_lcell_comb \Add1~48 (
// Equation(s):
// \Add1~48_combout  = ((dcifimemload_15 $ (\npc[26]~48_combout  $ (!\Add1~47 )))) # (GND)
// \Add1~49  = CARRY((dcifimemload_15 & ((\npc[26]~48_combout ) # (!\Add1~47 ))) # (!dcifimemload_15 & (\npc[26]~48_combout  & !\Add1~47 )))

	.dataa(dcifimemload_15),
	.datab(\npc[26]~48_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~47 ),
	.combout(\Add1~48_combout ),
	.cout(\Add1~49 ));
// synopsys translate_off
defparam \Add1~48 .lut_mask = 16'h698E;
defparam \Add1~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N20
cycloneive_lcell_comb \Add1~50 (
// Equation(s):
// \Add1~50_combout  = (dcifimemload_15 & ((\npc[27]~50_combout  & (\Add1~49  & VCC)) # (!\npc[27]~50_combout  & (!\Add1~49 )))) # (!dcifimemload_15 & ((\npc[27]~50_combout  & (!\Add1~49 )) # (!\npc[27]~50_combout  & ((\Add1~49 ) # (GND)))))
// \Add1~51  = CARRY((dcifimemload_15 & (!\npc[27]~50_combout  & !\Add1~49 )) # (!dcifimemload_15 & ((!\Add1~49 ) # (!\npc[27]~50_combout ))))

	.dataa(dcifimemload_15),
	.datab(\npc[27]~50_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~49 ),
	.combout(\Add1~50_combout ),
	.cout(\Add1~51 ));
// synopsys translate_off
defparam \Add1~50 .lut_mask = 16'h9617;
defparam \Add1~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N22
cycloneive_lcell_comb \Add1~52 (
// Equation(s):
// \Add1~52_combout  = ((dcifimemload_15 $ (\npc[28]~52_combout  $ (!\Add1~51 )))) # (GND)
// \Add1~53  = CARRY((dcifimemload_15 & ((\npc[28]~52_combout ) # (!\Add1~51 ))) # (!dcifimemload_15 & (\npc[28]~52_combout  & !\Add1~51 )))

	.dataa(dcifimemload_15),
	.datab(\npc[28]~52_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~51 ),
	.combout(\Add1~52_combout ),
	.cout(\Add1~53 ));
// synopsys translate_off
defparam \Add1~52 .lut_mask = 16'h698E;
defparam \Add1~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N24
cycloneive_lcell_comb \Add1~54 (
// Equation(s):
// \Add1~54_combout  = (dcifimemload_15 & ((\npc[29]~54_combout  & (\Add1~53  & VCC)) # (!\npc[29]~54_combout  & (!\Add1~53 )))) # (!dcifimemload_15 & ((\npc[29]~54_combout  & (!\Add1~53 )) # (!\npc[29]~54_combout  & ((\Add1~53 ) # (GND)))))
// \Add1~55  = CARRY((dcifimemload_15 & (!\npc[29]~54_combout  & !\Add1~53 )) # (!dcifimemload_15 & ((!\Add1~53 ) # (!\npc[29]~54_combout ))))

	.dataa(dcifimemload_15),
	.datab(\npc[29]~54_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~53 ),
	.combout(\Add1~54_combout ),
	.cout(\Add1~55 ));
// synopsys translate_off
defparam \Add1~54 .lut_mask = 16'h9617;
defparam \Add1~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N8
cycloneive_lcell_comb \PC[29]~1 (
// Equation(s):
// \PC[29]~1_combout  = (cuifPCSrc_1 & (Mux2)) # (!cuifPCSrc_1 & ((\Add1~54_combout )))

	.dataa(Mux2),
	.datab(cuifPCSrc_1),
	.datac(gnd),
	.datad(\Add1~54_combout ),
	.cin(gnd),
	.combout(\PC[29]~1_combout ),
	.cout());
// synopsys translate_off
defparam \PC[29]~1 .lut_mask = 16'hBB88;
defparam \PC[29]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N16
cycloneive_lcell_comb \PC[28]~0 (
// Equation(s):
// \PC[28]~0_combout  = (cuifPCSrc_1 & (Mux3)) # (!cuifPCSrc_1 & ((\Add1~52_combout )))

	.dataa(Mux3),
	.datab(cuifPCSrc_1),
	.datac(gnd),
	.datad(\Add1~52_combout ),
	.cin(gnd),
	.combout(\PC[28]~0_combout ),
	.cout());
// synopsys translate_off
defparam \PC[28]~0 .lut_mask = 16'hBB88;
defparam \PC[28]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N26
cycloneive_lcell_comb \npc[30]~56 (
// Equation(s):
// \npc[30]~56_combout  = (PC_30 & (\npc[29]~55  $ (GND))) # (!PC_30 & (!\npc[29]~55  & VCC))
// \npc[30]~57  = CARRY((PC_30 & !\npc[29]~55 ))

	.dataa(gnd),
	.datab(PC_30),
	.datac(gnd),
	.datad(vcc),
	.cin(\npc[29]~55 ),
	.combout(\npc[30]~56_combout ),
	.cout(\npc[30]~57 ));
// synopsys translate_off
defparam \npc[30]~56 .lut_mask = 16'hC30C;
defparam \npc[30]~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N28
cycloneive_lcell_comb \npc[31]~58 (
// Equation(s):
// \npc[31]~58_combout  = \npc[30]~57  $ (PC_31)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(PC_31),
	.cin(\npc[30]~57 ),
	.combout(\npc[31]~58_combout ),
	.cout());
// synopsys translate_off
defparam \npc[31]~58 .lut_mask = 16'h0FF0;
defparam \npc[31]~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N26
cycloneive_lcell_comb \Add1~56 (
// Equation(s):
// \Add1~56_combout  = ((\npc[30]~56_combout  $ (dcifimemload_15 $ (!\Add1~55 )))) # (GND)
// \Add1~57  = CARRY((\npc[30]~56_combout  & ((dcifimemload_15) # (!\Add1~55 ))) # (!\npc[30]~56_combout  & (dcifimemload_15 & !\Add1~55 )))

	.dataa(\npc[30]~56_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~55 ),
	.combout(\Add1~56_combout ),
	.cout(\Add1~57 ));
// synopsys translate_off
defparam \Add1~56 .lut_mask = 16'h698E;
defparam \Add1~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N28
cycloneive_lcell_comb \Add1~58 (
// Equation(s):
// \Add1~58_combout  = dcifimemload_15 $ (\Add1~57  $ (\npc[31]~58_combout ))

	.dataa(gnd),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(\npc[31]~58_combout ),
	.cin(\Add1~57 ),
	.combout(\Add1~58_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~58 .lut_mask = 16'hC33C;
defparam \Add1~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N28
cycloneive_lcell_comb \PC[31]~3 (
// Equation(s):
// \PC[31]~3_combout  = (cuifPCSrc_1 & (Mux0)) # (!cuifPCSrc_1 & ((\Add1~58_combout )))

	.dataa(cuifPCSrc_1),
	.datab(Mux0),
	.datac(gnd),
	.datad(\Add1~58_combout ),
	.cin(gnd),
	.combout(\PC[31]~3_combout ),
	.cout());
// synopsys translate_off
defparam \PC[31]~3 .lut_mask = 16'hDD88;
defparam \PC[31]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N30
cycloneive_lcell_comb \PC[30]~2 (
// Equation(s):
// \PC[30]~2_combout  = (cuifPCSrc_1 & (Mux1)) # (!cuifPCSrc_1 & ((\Add1~56_combout )))

	.dataa(cuifPCSrc_1),
	.datab(Mux1),
	.datac(gnd),
	.datad(\Add1~56_combout ),
	.cin(gnd),
	.combout(\PC[30]~2_combout ),
	.cout());
// synopsys translate_off
defparam \PC[30]~2 .lut_mask = 16'hDD88;
defparam \PC[30]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N26
cycloneive_lcell_comb \Mux30~2 (
// Equation(s):
// \Mux30~2_combout  = (!cuifPCSrc_0 & ((dcifimemload_25 & ((Mux30))) # (!dcifimemload_25 & (Mux301))))

	.dataa(dcifimemload_25),
	.datab(Mux301),
	.datac(Mux30),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~2 .lut_mask = 16'h00E4;
defparam \Mux30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N16
cycloneive_lcell_comb \PC[1]~4 (
// Equation(s):
// \PC[1]~4_combout  = (ccifiwait_0 & ((always0) # ((Equal31) # (Equal2))))

	.dataa(always0),
	.datab(\pcuif.ihit ),
	.datac(Equal3),
	.datad(Equal2),
	.cin(gnd),
	.combout(\PC[1]~4_combout ),
	.cout());
// synopsys translate_off
defparam \PC[1]~4 .lut_mask = 16'hCCC8;
defparam \PC[1]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N4
cycloneive_lcell_comb \Mux31~2 (
// Equation(s):
// \Mux31~2_combout  = (!cuifPCSrc_0 & ((dcifimemload_25 & (Mux31)) # (!dcifimemload_25 & ((Mux311)))))

	.dataa(Mux31),
	.datab(dcifimemload_25),
	.datac(cuifPCSrc_0),
	.datad(Mux311),
	.cin(gnd),
	.combout(\Mux31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~2 .lut_mask = 16'h0B08;
defparam \Mux31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N24
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (cuifPCSrc_1 & (((!cuifPCSrc_0)))) # (!cuifPCSrc_1 & ((cuifPCSrc_0 & ((\npc[3]~2_combout ))) # (!cuifPCSrc_0 & (\Add1~2_combout ))))

	.dataa(\Add1~2_combout ),
	.datab(cuifPCSrc_1),
	.datac(\npc[3]~2_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'h30EE;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N0
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (cuifPCSrc_1 & ((\Mux28~0_combout  & (Mux28)) # (!\Mux28~0_combout  & ((dcifimemload_1))))) # (!cuifPCSrc_1 & (((\Mux28~0_combout ))))

	.dataa(Mux28),
	.datab(cuifPCSrc_1),
	.datac(dcifimemload_1),
	.datad(\Mux28~0_combout ),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hBBC0;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N14
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (cuifPCSrc_1 & (((dcifimemload_0) # (!cuifPCSrc_0)))) # (!cuifPCSrc_1 & (\npc[2]~0_combout  & ((cuifPCSrc_0))))

	.dataa(\npc[2]~0_combout ),
	.datab(cuifPCSrc_1),
	.datac(dcifimemload_0),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hE2CC;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N2
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// \Mux29~1_combout  = (\Mux29~0_combout  & ((Mux292) # ((cuifPCSrc_0)))) # (!\Mux29~0_combout  & (((\Add1~0_combout  & !cuifPCSrc_0))))

	.dataa(Mux29),
	.datab(\Add1~0_combout ),
	.datac(\Mux29~0_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hF0AC;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N26
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (cuifPCSrc_1 & (((!cuifPCSrc_0)))) # (!cuifPCSrc_1 & ((cuifPCSrc_0 & (\npc[5]~6_combout )) # (!cuifPCSrc_0 & ((\Add1~6_combout )))))

	.dataa(\npc[5]~6_combout ),
	.datab(\Add1~6_combout ),
	.datac(cuifPCSrc_1),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'h0AFC;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N12
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (cuifPCSrc_1 & ((\Mux26~0_combout  & ((Mux26))) # (!\Mux26~0_combout  & (dcifimemload_3)))) # (!cuifPCSrc_1 & (((\Mux26~0_combout ))))

	.dataa(dcifimemload_3),
	.datab(cuifPCSrc_1),
	.datac(\Mux26~0_combout ),
	.datad(Mux26),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hF838;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N4
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (cuifPCSrc_1 & (((dcifimemload_2) # (!cuifPCSrc_0)))) # (!cuifPCSrc_1 & (\npc[4]~4_combout  & ((cuifPCSrc_0))))

	.dataa(\npc[4]~4_combout ),
	.datab(cuifPCSrc_1),
	.datac(dcifimemload_2),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hE2CC;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N2
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// \Mux27~1_combout  = (\Mux27~0_combout  & ((Mux272) # ((cuifPCSrc_0)))) # (!\Mux27~0_combout  & (((\Add1~4_combout  & !cuifPCSrc_0))))

	.dataa(Mux27),
	.datab(\Add1~4_combout ),
	.datac(\Mux27~0_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hF0AC;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N22
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (cuifPCSrc_1 & (((!cuifPCSrc_0)))) # (!cuifPCSrc_1 & ((cuifPCSrc_0 & ((\npc[7]~10_combout ))) # (!cuifPCSrc_0 & (\Add1~10_combout ))))

	.dataa(cuifPCSrc_1),
	.datab(\Add1~10_combout ),
	.datac(\npc[7]~10_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'h50EE;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N0
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// \Mux24~1_combout  = (cuifPCSrc_1 & ((\Mux24~0_combout  & (Mux242)) # (!\Mux24~0_combout  & ((dcifimemload_5))))) # (!cuifPCSrc_1 & (((\Mux24~0_combout ))))

	.dataa(cuifPCSrc_1),
	.datab(Mux24),
	.datac(\Mux24~0_combout ),
	.datad(dcifimemload_5),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hDAD0;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N24
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (cuifPCSrc_1 & ((dcifimemload_4) # ((!cuifPCSrc_0)))) # (!cuifPCSrc_1 & (((\npc[6]~8_combout  & cuifPCSrc_0))))

	.dataa(cuifPCSrc_1),
	.datab(dcifimemload_4),
	.datac(\npc[6]~8_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hD8AA;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N4
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (cuifPCSrc_0 & (((\Mux25~0_combout )))) # (!cuifPCSrc_0 & ((\Mux25~0_combout  & (Mux252)) # (!\Mux25~0_combout  & ((\Add1~8_combout )))))

	.dataa(Mux25),
	.datab(cuifPCSrc_0),
	.datac(\Add1~8_combout ),
	.datad(\Mux25~0_combout ),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hEE30;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N2
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (cuifPCSrc_1 & (((!cuifPCSrc_0)))) # (!cuifPCSrc_1 & ((cuifPCSrc_0 & (\npc[9]~14_combout )) # (!cuifPCSrc_0 & ((\Add1~14_combout )))))

	.dataa(cuifPCSrc_1),
	.datab(\npc[9]~14_combout ),
	.datac(\Add1~14_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'h44FA;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N30
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// \Mux22~1_combout  = (cuifPCSrc_1 & ((\Mux22~0_combout  & ((Mux22))) # (!\Mux22~0_combout  & (dcifimemload_7)))) # (!cuifPCSrc_1 & (((\Mux22~0_combout ))))

	.dataa(cuifPCSrc_1),
	.datab(dcifimemload_7),
	.datac(Mux22),
	.datad(\Mux22~0_combout ),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'hF588;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N28
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (cuifPCSrc_0 & ((cuifPCSrc_1 & (dcifimemload_6)) # (!cuifPCSrc_1 & ((\npc[8]~12_combout ))))) # (!cuifPCSrc_0 & (((cuifPCSrc_1))))

	.dataa(dcifimemload_6),
	.datab(\npc[8]~12_combout ),
	.datac(cuifPCSrc_0),
	.datad(cuifPCSrc_1),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hAFC0;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N8
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// \Mux23~1_combout  = (cuifPCSrc_0 & (((\Mux23~0_combout )))) # (!cuifPCSrc_0 & ((\Mux23~0_combout  & ((Mux23))) # (!\Mux23~0_combout  & (\Add1~12_combout ))))

	.dataa(\Add1~12_combout ),
	.datab(Mux23),
	.datac(cuifPCSrc_0),
	.datad(\Mux23~0_combout ),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'hFC0A;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N2
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (cuifPCSrc_1 & (((!cuifPCSrc_0)))) # (!cuifPCSrc_1 & ((cuifPCSrc_0 & ((\npc[11]~18_combout ))) # (!cuifPCSrc_0 & (\Add1~18_combout ))))

	.dataa(cuifPCSrc_1),
	.datab(\Add1~18_combout ),
	.datac(\npc[11]~18_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'h50EE;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N12
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// \Mux20~1_combout  = (cuifPCSrc_1 & ((\Mux20~0_combout  & (Mux20)) # (!\Mux20~0_combout  & ((dcifimemload_9))))) # (!cuifPCSrc_1 & (((\Mux20~0_combout ))))

	.dataa(Mux20),
	.datab(dcifimemload_9),
	.datac(cuifPCSrc_1),
	.datad(\Mux20~0_combout ),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'hAFC0;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N10
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (cuifPCSrc_0 & ((cuifPCSrc_1 & (dcifimemload_8)) # (!cuifPCSrc_1 & ((\npc[10]~16_combout ))))) # (!cuifPCSrc_0 & (((cuifPCSrc_1))))

	.dataa(dcifimemload_8),
	.datab(\npc[10]~16_combout ),
	.datac(cuifPCSrc_0),
	.datad(cuifPCSrc_1),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hAFC0;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N30
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// \Mux21~1_combout  = (cuifPCSrc_0 & (((\Mux21~0_combout )))) # (!cuifPCSrc_0 & ((\Mux21~0_combout  & ((Mux21))) # (!\Mux21~0_combout  & (\Add1~16_combout ))))

	.dataa(\Add1~16_combout ),
	.datab(Mux21),
	.datac(cuifPCSrc_0),
	.datad(\Mux21~0_combout ),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'hFC0A;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N16
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (cuifPCSrc_1 & (((!cuifPCSrc_0)))) # (!cuifPCSrc_1 & ((cuifPCSrc_0 & (\npc[13]~22_combout )) # (!cuifPCSrc_0 & ((\Add1~22_combout )))))

	.dataa(\npc[13]~22_combout ),
	.datab(cuifPCSrc_1),
	.datac(cuifPCSrc_0),
	.datad(\Add1~22_combout ),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'h2F2C;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N4
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// \Mux18~1_combout  = (cuifPCSrc_1 & ((\Mux18~0_combout  & (Mux18)) # (!\Mux18~0_combout  & ((dcifimemload_11))))) # (!cuifPCSrc_1 & (((\Mux18~0_combout ))))

	.dataa(Mux18),
	.datab(cuifPCSrc_1),
	.datac(dcifimemload_11),
	.datad(\Mux18~0_combout ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'hBBC0;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N6
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (cuifPCSrc_1 & ((dcifimemload_10) # ((!cuifPCSrc_0)))) # (!cuifPCSrc_1 & (((cuifPCSrc_0 & \npc[12]~20_combout ))))

	.dataa(dcifimemload_10),
	.datab(cuifPCSrc_1),
	.datac(cuifPCSrc_0),
	.datad(\npc[12]~20_combout ),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'hBC8C;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N22
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// \Mux19~1_combout  = (cuifPCSrc_0 & (((\Mux19~0_combout )))) # (!cuifPCSrc_0 & ((\Mux19~0_combout  & (Mux19)) # (!\Mux19~0_combout  & ((\Add1~20_combout )))))

	.dataa(Mux19),
	.datab(\Add1~20_combout ),
	.datac(cuifPCSrc_0),
	.datad(\Mux19~0_combout ),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hFA0C;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N24
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (cuifPCSrc_1 & (((!cuifPCSrc_0)))) # (!cuifPCSrc_1 & ((cuifPCSrc_0 & (\npc[15]~26_combout )) # (!cuifPCSrc_0 & ((\Add1~26_combout )))))

	.dataa(\npc[15]~26_combout ),
	.datab(cuifPCSrc_1),
	.datac(cuifPCSrc_0),
	.datad(\Add1~26_combout ),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'h2F2C;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N20
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// \Mux16~1_combout  = (cuifPCSrc_1 & ((\Mux16~0_combout  & ((Mux16))) # (!\Mux16~0_combout  & (dcifimemload_13)))) # (!cuifPCSrc_1 & (((\Mux16~0_combout ))))

	.dataa(dcifimemload_13),
	.datab(cuifPCSrc_1),
	.datac(Mux16),
	.datad(\Mux16~0_combout ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hF388;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N18
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (cuifPCSrc_0 & ((cuifPCSrc_1 & (dcifimemload_12)) # (!cuifPCSrc_1 & ((\npc[14]~24_combout ))))) # (!cuifPCSrc_0 & (((cuifPCSrc_1))))

	.dataa(dcifimemload_12),
	.datab(\npc[14]~24_combout ),
	.datac(cuifPCSrc_0),
	.datad(cuifPCSrc_1),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hAFC0;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N14
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// \Mux17~1_combout  = (cuifPCSrc_0 & (((\Mux17~0_combout )))) # (!cuifPCSrc_0 & ((\Mux17~0_combout  & (Mux17)) # (!\Mux17~0_combout  & ((\Add1~24_combout )))))

	.dataa(Mux17),
	.datab(\Add1~24_combout ),
	.datac(cuifPCSrc_0),
	.datad(\Mux17~0_combout ),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hFA0C;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N12
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (cuifPCSrc_0 & (((\npc[17]~30_combout  & !cuifPCSrc_1)))) # (!cuifPCSrc_0 & ((\Add1~30_combout ) # ((cuifPCSrc_1))))

	.dataa(\Add1~30_combout ),
	.datab(\npc[17]~30_combout ),
	.datac(cuifPCSrc_0),
	.datad(cuifPCSrc_1),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'h0FCA;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N0
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// \Mux14~1_combout  = (\Mux14~0_combout  & (((Mux14)) # (!cuifPCSrc_1))) # (!\Mux14~0_combout  & (cuifPCSrc_1 & (dcifimemload_15)))

	.dataa(\Mux14~0_combout ),
	.datab(cuifPCSrc_1),
	.datac(dcifimemload_15),
	.datad(Mux14),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hEA62;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N26
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (cuifPCSrc_1 & ((dcifimemload_14) # ((!cuifPCSrc_0)))) # (!cuifPCSrc_1 & (((\npc[16]~28_combout  & cuifPCSrc_0))))

	.dataa(cuifPCSrc_1),
	.datab(dcifimemload_14),
	.datac(\npc[16]~28_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hD8AA;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N0
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// \Mux15~1_combout  = (\Mux15~0_combout  & ((Mux15) # ((cuifPCSrc_0)))) # (!\Mux15~0_combout  & (((\Add1~28_combout  & !cuifPCSrc_0))))

	.dataa(Mux15),
	.datab(\Add1~28_combout ),
	.datac(\Mux15~0_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hF0AC;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N12
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (cuifPCSrc_1 & (((!cuifPCSrc_0)))) # (!cuifPCSrc_1 & ((cuifPCSrc_0 & (\npc[19]~34_combout )) # (!cuifPCSrc_0 & ((\Add1~34_combout )))))

	.dataa(cuifPCSrc_1),
	.datab(\npc[19]~34_combout ),
	.datac(\Add1~34_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'h44FA;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N10
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// \Mux12~1_combout  = (cuifPCSrc_1 & ((\Mux12~0_combout  & (Mux12)) # (!\Mux12~0_combout  & ((dcifimemload_17))))) # (!cuifPCSrc_1 & (((\Mux12~0_combout ))))

	.dataa(cuifPCSrc_1),
	.datab(Mux12),
	.datac(dcifimemload_17),
	.datad(\Mux12~0_combout ),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hDDA0;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N22
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (cuifPCSrc_1 & (((dcifimemload_16) # (!cuifPCSrc_0)))) # (!cuifPCSrc_1 & (\npc[18]~32_combout  & ((cuifPCSrc_0))))

	.dataa(cuifPCSrc_1),
	.datab(\npc[18]~32_combout ),
	.datac(dcifimemload_16),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hE4AA;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N28
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// \Mux13~1_combout  = (\Mux13~0_combout  & ((Mux13) # ((cuifPCSrc_0)))) # (!\Mux13~0_combout  & (((\Add1~32_combout  & !cuifPCSrc_0))))

	.dataa(Mux13),
	.datab(\Add1~32_combout ),
	.datac(\Mux13~0_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hF0AC;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N24
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (cuifPCSrc_0 & (\npc[21]~38_combout  & ((!cuifPCSrc_1)))) # (!cuifPCSrc_0 & (((\Add1~38_combout ) # (cuifPCSrc_1))))

	.dataa(\npc[21]~38_combout ),
	.datab(\Add1~38_combout ),
	.datac(cuifPCSrc_0),
	.datad(cuifPCSrc_1),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'h0FAC;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N20
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// \Mux10~1_combout  = (cuifPCSrc_1 & ((\Mux10~0_combout  & (Mux10)) # (!\Mux10~0_combout  & ((dcifimemload_19))))) # (!cuifPCSrc_1 & (((\Mux10~0_combout ))))

	.dataa(Mux10),
	.datab(dcifimemload_19),
	.datac(cuifPCSrc_1),
	.datad(\Mux10~0_combout ),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hAFC0;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N4
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (cuifPCSrc_1 & (((dcifimemload_18) # (!cuifPCSrc_0)))) # (!cuifPCSrc_1 & (\npc[20]~36_combout  & ((cuifPCSrc_0))))

	.dataa(cuifPCSrc_1),
	.datab(\npc[20]~36_combout ),
	.datac(dcifimemload_18),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hE4AA;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N2
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// \Mux11~1_combout  = (\Mux11~0_combout  & ((Mux11) # ((cuifPCSrc_0)))) # (!\Mux11~0_combout  & (((\Add1~36_combout  & !cuifPCSrc_0))))

	.dataa(Mux11),
	.datab(\Add1~36_combout ),
	.datac(\Mux11~0_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hF0AC;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N16
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (cuifPCSrc_1 & (((!cuifPCSrc_0)))) # (!cuifPCSrc_1 & ((cuifPCSrc_0 & (\npc[23]~42_combout )) # (!cuifPCSrc_0 & ((\Add1~42_combout )))))

	.dataa(\npc[23]~42_combout ),
	.datab(cuifPCSrc_1),
	.datac(\Add1~42_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'h22FC;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N4
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// \Mux8~1_combout  = (cuifPCSrc_1 & ((\Mux8~0_combout  & (Mux8)) # (!\Mux8~0_combout  & ((dcifimemload_21))))) # (!cuifPCSrc_1 & (((\Mux8~0_combout ))))

	.dataa(Mux8),
	.datab(cuifPCSrc_1),
	.datac(dcifimemload_21),
	.datad(\Mux8~0_combout ),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hBBC0;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N6
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (cuifPCSrc_1 & (((dcifimemload_20) # (!cuifPCSrc_0)))) # (!cuifPCSrc_1 & (\npc[22]~40_combout  & ((cuifPCSrc_0))))

	.dataa(cuifPCSrc_1),
	.datab(\npc[22]~40_combout ),
	.datac(dcifimemload_20),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hE4AA;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N16
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// \Mux9~1_combout  = (cuifPCSrc_0 & (((\Mux9~0_combout )))) # (!cuifPCSrc_0 & ((\Mux9~0_combout  & (Mux9)) # (!\Mux9~0_combout  & ((\Add1~40_combout )))))

	.dataa(Mux9),
	.datab(cuifPCSrc_0),
	.datac(\Add1~40_combout ),
	.datad(\Mux9~0_combout ),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hEE30;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N10
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (cuifPCSrc_1 & (((!cuifPCSrc_0)))) # (!cuifPCSrc_1 & ((cuifPCSrc_0 & (\npc[25]~46_combout )) # (!cuifPCSrc_0 & ((\Add1~46_combout )))))

	.dataa(\npc[25]~46_combout ),
	.datab(\Add1~46_combout ),
	.datac(cuifPCSrc_1),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'h0AFC;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N8
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// \Mux6~1_combout  = (cuifPCSrc_1 & ((\Mux6~0_combout  & (Mux6)) # (!\Mux6~0_combout  & ((dcifimemload_23))))) # (!cuifPCSrc_1 & (((\Mux6~0_combout ))))

	.dataa(Mux6),
	.datab(dcifimemload_23),
	.datac(cuifPCSrc_1),
	.datad(\Mux6~0_combout ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hAFC0;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N8
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (cuifPCSrc_1 & (((dcifimemload_22) # (!cuifPCSrc_0)))) # (!cuifPCSrc_1 & (\npc[24]~44_combout  & ((cuifPCSrc_0))))

	.dataa(\npc[24]~44_combout ),
	.datab(cuifPCSrc_1),
	.datac(dcifimemload_22),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hE2CC;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N30
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// \Mux7~1_combout  = (\Mux7~0_combout  & (((Mux72) # (cuifPCSrc_0)))) # (!\Mux7~0_combout  & (\Add1~44_combout  & ((!cuifPCSrc_0))))

	.dataa(\Add1~44_combout ),
	.datab(Mux7),
	.datac(\Mux7~0_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hF0CA;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N28
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (cuifPCSrc_1 & (((!cuifPCSrc_0)))) # (!cuifPCSrc_1 & ((cuifPCSrc_0 & ((\npc[27]~50_combout ))) # (!cuifPCSrc_0 & (\Add1~50_combout ))))

	.dataa(cuifPCSrc_1),
	.datab(\Add1~50_combout ),
	.datac(\npc[27]~50_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'h50EE;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N12
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// \Mux4~1_combout  = (cuifPCSrc_1 & ((\Mux4~0_combout  & ((Mux4))) # (!\Mux4~0_combout  & (dcifimemload_25)))) # (!cuifPCSrc_1 & (((\Mux4~0_combout ))))

	.dataa(dcifimemload_25),
	.datab(Mux4),
	.datac(cuifPCSrc_1),
	.datad(\Mux4~0_combout ),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hCFA0;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N14
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = (cuifPCSrc_1 & (((dcifimemload_24) # (!cuifPCSrc_0)))) # (!cuifPCSrc_1 & (\npc[26]~48_combout  & ((cuifPCSrc_0))))

	.dataa(cuifPCSrc_1),
	.datab(\npc[26]~48_combout ),
	.datac(dcifimemload_24),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hE4AA;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N24
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// \Mux5~1_combout  = (\Mux5~0_combout  & (((Mux5) # (cuifPCSrc_0)))) # (!\Mux5~0_combout  & (\Add1~48_combout  & ((!cuifPCSrc_0))))

	.dataa(\Add1~48_combout ),
	.datab(Mux5),
	.datac(\Mux5~0_combout ),
	.datad(cuifPCSrc_0),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'hF0CA;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module register_file (
	ramiframload_16,
	ramiframload_17,
	ccifiwait_0,
	dcifimemload_19,
	dcifimemload_18,
	instr_16,
	dcifimemload_16,
	instr_17,
	dcifimemload_17,
	Mux63,
	Mux631,
	dcifimemload_24,
	dcifimemload_23,
	dcifimemload_21,
	dcifimemload_22,
	Mux30,
	Mux301,
	dcifimemload_25,
	Mux302,
	Mux0,
	Mux32,
	Mux321,
	Mux1,
	Mux33,
	Mux331,
	Mux2,
	Mux34,
	Mux341,
	Mux3,
	Mux35,
	Mux351,
	Mux4,
	Mux36,
	Mux361,
	Mux5,
	Mux37,
	Mux371,
	Mux6,
	Mux38,
	Mux381,
	Mux7,
	Mux71,
	Mux72,
	Mux39,
	Mux391,
	Mux8,
	Mux40,
	Mux401,
	Mux9,
	Mux41,
	Mux411,
	Mux10,
	Mux42,
	Mux421,
	Mux11,
	Mux43,
	Mux431,
	Mux12,
	Mux44,
	Mux441,
	Mux13,
	Mux45,
	Mux451,
	Mux14,
	Mux46,
	Mux461,
	Mux15,
	Mux47,
	Mux471,
	Mux16,
	Mux48,
	Mux481,
	Mux17,
	Mux49,
	Mux491,
	Mux18,
	Mux50,
	Mux501,
	Mux19,
	Mux51,
	Mux511,
	Mux20,
	Mux52,
	Mux521,
	Mux21,
	Mux53,
	Mux531,
	Mux22,
	Mux54,
	Mux541,
	Mux23,
	Mux55,
	Mux551,
	Mux24,
	Mux241,
	Mux242,
	Mux56,
	Mux561,
	Mux25,
	Mux251,
	Mux252,
	Mux57,
	Mux571,
	Mux26,
	Mux58,
	Mux581,
	Mux27,
	Mux271,
	Mux272,
	Mux59,
	Mux591,
	Mux28,
	Mux60,
	Mux601,
	Mux29,
	Mux291,
	Mux292,
	Mux61,
	Mux611,
	Mux62,
	Mux621,
	Mux31,
	Mux311,
	Mux312,
	wdat,
	cuifRegWEN,
	wsel,
	wsel1,
	wsel2,
	wsel3,
	wsel4,
	wdat1,
	wdat2,
	wdat3,
	wdat4,
	wdat5,
	wdat6,
	wdat7,
	wdat8,
	wdat9,
	wdat10,
	wdat11,
	wdat12,
	wdat13,
	wdat14,
	wdat15,
	wdat16,
	wdat17,
	wdat18,
	wdat19,
	wdat20,
	wdat21,
	wdat22,
	wdat23,
	wdat24,
	wdat25,
	wdat26,
	wdat27,
	wdat28,
	wdat29,
	wdat30,
	wdat31,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	ramiframload_16;
input 	ramiframload_17;
input 	ccifiwait_0;
input 	dcifimemload_19;
input 	dcifimemload_18;
input 	instr_16;
input 	dcifimemload_16;
input 	instr_17;
input 	dcifimemload_17;
output 	Mux63;
output 	Mux631;
input 	dcifimemload_24;
input 	dcifimemload_23;
input 	dcifimemload_21;
input 	dcifimemload_22;
output 	Mux30;
output 	Mux301;
input 	dcifimemload_25;
output 	Mux302;
output 	Mux0;
output 	Mux32;
output 	Mux321;
output 	Mux1;
output 	Mux33;
output 	Mux331;
output 	Mux2;
output 	Mux34;
output 	Mux341;
output 	Mux3;
output 	Mux35;
output 	Mux351;
output 	Mux4;
output 	Mux36;
output 	Mux361;
output 	Mux5;
output 	Mux37;
output 	Mux371;
output 	Mux6;
output 	Mux38;
output 	Mux381;
output 	Mux7;
output 	Mux71;
output 	Mux72;
output 	Mux39;
output 	Mux391;
output 	Mux8;
output 	Mux40;
output 	Mux401;
output 	Mux9;
output 	Mux41;
output 	Mux411;
output 	Mux10;
output 	Mux42;
output 	Mux421;
output 	Mux11;
output 	Mux43;
output 	Mux431;
output 	Mux12;
output 	Mux44;
output 	Mux441;
output 	Mux13;
output 	Mux45;
output 	Mux451;
output 	Mux14;
output 	Mux46;
output 	Mux461;
output 	Mux15;
output 	Mux47;
output 	Mux471;
output 	Mux16;
output 	Mux48;
output 	Mux481;
output 	Mux17;
output 	Mux49;
output 	Mux491;
output 	Mux18;
output 	Mux50;
output 	Mux501;
output 	Mux19;
output 	Mux51;
output 	Mux511;
output 	Mux20;
output 	Mux52;
output 	Mux521;
output 	Mux21;
output 	Mux53;
output 	Mux531;
output 	Mux22;
output 	Mux54;
output 	Mux541;
output 	Mux23;
output 	Mux55;
output 	Mux551;
output 	Mux24;
output 	Mux241;
output 	Mux242;
output 	Mux56;
output 	Mux561;
output 	Mux25;
output 	Mux251;
output 	Mux252;
output 	Mux57;
output 	Mux571;
output 	Mux26;
output 	Mux58;
output 	Mux581;
output 	Mux27;
output 	Mux271;
output 	Mux272;
output 	Mux59;
output 	Mux591;
output 	Mux28;
output 	Mux60;
output 	Mux601;
output 	Mux29;
output 	Mux291;
output 	Mux292;
output 	Mux61;
output 	Mux611;
output 	Mux62;
output 	Mux621;
output 	Mux31;
output 	Mux311;
output 	Mux312;
input 	wdat;
input 	cuifRegWEN;
input 	wsel;
input 	wsel1;
input 	wsel2;
input 	wsel3;
input 	wsel4;
input 	wdat1;
input 	wdat2;
input 	wdat3;
input 	wdat4;
input 	wdat5;
input 	wdat6;
input 	wdat7;
input 	wdat8;
input 	wdat9;
input 	wdat10;
input 	wdat11;
input 	wdat12;
input 	wdat13;
input 	wdat14;
input 	wdat15;
input 	wdat16;
input 	wdat17;
input 	wdat18;
input 	wdat19;
input 	wdat20;
input 	wdat21;
input 	wdat22;
input 	wdat23;
input 	wdat24;
input 	wdat25;
input 	wdat26;
input 	wdat27;
input 	wdat28;
input 	wdat29;
input 	wdat30;
input 	wdat31;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \my_reg[4][0]~q ;
wire \Mux63~12_combout ;
wire \Mux63~16_combout ;
wire \my_reg[22][1]~q ;
wire \my_reg[24][1]~q ;
wire \Mux0~4_combout ;
wire \my_reg[10][31]~q ;
wire \my_reg[5][31]~q ;
wire \Mux32~2_combout ;
wire \my_reg[10][30]~q ;
wire \my_reg[17][29]~q ;
wire \my_reg[21][28]~q ;
wire \my_reg[12][28]~q ;
wire \Mux3~17_combout ;
wire \Mux5~4_combout ;
wire \my_reg[23][26]~q ;
wire \my_reg[2][26]~q ;
wire \my_reg[1][25]~q ;
wire \Mux6~14_combout ;
wire \Mux8~10_combout ;
wire \my_reg[13][23]~q ;
wire \my_reg[5][22]~q ;
wire \my_reg[3][22]~q ;
wire \Mux41~2_combout ;
wire \Mux41~4_combout ;
wire \my_reg[1][21]~q ;
wire \Mux10~14_combout ;
wire \my_reg[12][21]~q ;
wire \Mux10~17_combout ;
wire \Mux42~2_combout ;
wire \Mux11~12_combout ;
wire \Mux11~13_combout ;
wire \my_reg[27][19]~q ;
wire \my_reg[5][18]~q ;
wire \Mux45~2_combout ;
wire \my_reg[20][17]~q ;
wire \Mux15~2_combout ;
wire \my_reg[30][16]~q ;
wire \Mux15~3_combout ;
wire \my_reg[20][15]~q ;
wire \my_reg[27][15]~q ;
wire \Mux48~14_combout ;
wire \my_reg[17][14]~q ;
wire \Mux17~0_combout ;
wire \my_reg[24][14]~q ;
wire \my_reg[5][14]~q ;
wire \Mux49~14_combout ;
wire \my_reg[18][13]~q ;
wire \Mux18~2_combout ;
wire \my_reg[30][13]~q ;
wire \Mux18~3_combout ;
wire \my_reg[1][13]~q ;
wire \Mux18~14_combout ;
wire \my_reg[12][13]~q ;
wire \my_reg[17][12]~q ;
wire \my_reg[22][12]~q ;
wire \my_reg[23][12]~q ;
wire \my_reg[5][12]~q ;
wire \Mux52~4_combout ;
wire \my_reg[17][10]~q ;
wire \Mux21~0_combout ;
wire \my_reg[17][9]~q ;
wire \Mux22~0_combout ;
wire \my_reg[30][9]~q ;
wire \my_reg[9][9]~q ;
wire \my_reg[21][8]~q ;
wire \my_reg[22][8]~q ;
wire \my_reg[24][7]~q ;
wire \my_reg[19][7]~q ;
wire \my_reg[17][6]~q ;
wire \my_reg[1][6]~q ;
wire \my_reg[25][5]~q ;
wire \my_reg[26][5]~q ;
wire \my_reg[24][3]~q ;
wire \my_reg[16][3]~q ;
wire \Mux28~4_combout ;
wire \Mux28~5_combout ;
wire \my_reg[20][2]~q ;
wire \my_reg[10][2]~q ;
wire \Mux62~14_combout ;
wire \Decoder0~50_combout ;
wire \my_reg[24][1]~feeder_combout ;
wire \my_reg[22][1]~feeder_combout ;
wire \my_reg[5][31]~feeder_combout ;
wire \my_reg[10][30]~feeder_combout ;
wire \my_reg[17][29]~feeder_combout ;
wire \my_reg[21][28]~feeder_combout ;
wire \my_reg[23][26]~feeder_combout ;
wire \my_reg[2][26]~feeder_combout ;
wire \my_reg[13][23]~feeder_combout ;
wire \my_reg[27][19]~feeder_combout ;
wire \my_reg[20][17]~feeder_combout ;
wire \my_reg[30][16]~feeder_combout ;
wire \my_reg[27][15]~feeder_combout ;
wire \my_reg[17][14]~feeder_combout ;
wire \my_reg[5][14]~feeder_combout ;
wire \my_reg[1][13]~feeder_combout ;
wire \my_reg[12][13]~feeder_combout ;
wire \my_reg[30][13]~feeder_combout ;
wire \my_reg[18][13]~feeder_combout ;
wire \my_reg[5][12]~feeder_combout ;
wire \my_reg[22][12]~feeder_combout ;
wire \my_reg[17][12]~feeder_combout ;
wire \my_reg[23][12]~feeder_combout ;
wire \my_reg[9][9]~feeder_combout ;
wire \my_reg[17][9]~feeder_combout ;
wire \my_reg[30][9]~feeder_combout ;
wire \my_reg[21][8]~feeder_combout ;
wire \my_reg[22][8]~feeder_combout ;
wire \my_reg[24][7]~feeder_combout ;
wire \my_reg[19][7]~feeder_combout ;
wire \my_reg[1][6]~feeder_combout ;
wire \my_reg[17][6]~feeder_combout ;
wire \my_reg[25][5]~feeder_combout ;
wire \my_reg[26][5]~feeder_combout ;
wire \my_reg[24][3]~feeder_combout ;
wire \my_reg[16][3]~feeder_combout ;
wire \my_reg[20][2]~feeder_combout ;
wire \my_reg[10][2]~feeder_combout ;
wire \Decoder0~15_combout ;
wire \Decoder0~16_combout ;
wire \my_reg[29][0]~q ;
wire \my_reg[25][0]~feeder_combout ;
wire \Decoder0~10_combout ;
wire \Decoder0~11_combout ;
wire \my_reg[25][0]~q ;
wire \my_reg[21][0]~feeder_combout ;
wire \Decoder0~12_combout ;
wire \Decoder0~13_combout ;
wire \my_reg[21][0]~q ;
wire \Mux63~0_combout ;
wire \Mux63~1_combout ;
wire \Decoder0~19_combout ;
wire \Decoder0~22_combout ;
wire \my_reg[30][0]~q ;
wire \Decoder0~17_combout ;
wire \Decoder0~21_combout ;
wire \my_reg[18][0]~q ;
wire \Decoder0~20_combout ;
wire \my_reg[26][0]~q ;
wire \Mux63~2_combout ;
wire \Mux63~3_combout ;
wire \Decoder0~24_combout ;
wire \my_reg[16][0]~q ;
wire \Decoder0~23_combout ;
wire \my_reg[20][0]~q ;
wire \Decoder0~26_combout ;
wire \my_reg[24][0]~q ;
wire \Mux63~4_combout ;
wire \Mux63~5_combout ;
wire \Mux63~6_combout ;
wire \Decoder0~30_combout ;
wire \my_reg[31][0]~q ;
wire \my_reg[27][0]~feeder_combout ;
wire \Decoder0~27_combout ;
wire \my_reg[27][0]~q ;
wire \my_reg[23][0]~feeder_combout ;
wire \Decoder0~28_combout ;
wire \my_reg[23][0]~q ;
wire \Mux63~7_combout ;
wire \Mux63~8_combout ;
wire \Decoder0~51_combout ;
wire \Decoder0~42_combout ;
wire \my_reg[2][0]~q ;
wire \Decoder0~41_combout ;
wire \my_reg[3][0]~q ;
wire \Decoder0~52_combout ;
wire \my_reg[1][0]~q ;
wire \Mux63~17_combout ;
wire \Mux63~18_combout ;
wire \Mux63~19_combout ;
wire \Decoder0~36_combout ;
wire \my_reg[6][0]~q ;
wire \Decoder0~40_combout ;
wire \my_reg[7][0]~q ;
wire \Decoder0~35_combout ;
wire \Decoder0~37_combout ;
wire \Decoder0~38_combout ;
wire \my_reg[5][0]~q ;
wire \Mux63~13_combout ;
wire \Mux63~14_combout ;
wire \Mux63~15_combout ;
wire \Mux63~20_combout ;
wire \my_reg[14][0]~feeder_combout ;
wire \Decoder0~49_combout ;
wire \Decoder0~43_combout ;
wire \my_reg[14][0]~q ;
wire \Decoder0~47_combout ;
wire \my_reg[15][0]~q ;
wire \my_reg[12][0]~feeder_combout ;
wire \Decoder0~31_combout ;
wire \Decoder0~44_combout ;
wire \Decoder0~46_combout ;
wire \my_reg[12][0]~q ;
wire \Decoder0~45_combout ;
wire \my_reg[13][0]~q ;
wire \Mux63~21_combout ;
wire \Mux63~22_combout ;
wire \Decoder0~34_combout ;
wire \my_reg[11][0]~q ;
wire \my_reg[10][0]~feeder_combout ;
wire \Decoder0~32_combout ;
wire \my_reg[10][0]~q ;
wire \Mux63~10_combout ;
wire \Decoder0~48_combout ;
wire \my_reg[9][0]~q ;
wire \Mux63~11_combout ;
wire \my_reg[25][1]~q ;
wire \my_reg[29][1]~feeder_combout ;
wire \my_reg[29][1]~q ;
wire \my_reg[21][1]~q ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \my_reg[20][1]~feeder_combout ;
wire \my_reg[20][1]~q ;
wire \my_reg[16][1]~q ;
wire \Mux30~4_combout ;
wire \Mux30~5_combout ;
wire \my_reg[30][1]~q ;
wire \my_reg[18][1]~q ;
wire \Mux30~2_combout ;
wire \Mux30~3_combout ;
wire \Mux30~6_combout ;
wire \my_reg[27][1]~feeder_combout ;
wire \my_reg[27][1]~q ;
wire \my_reg[31][1]~q ;
wire \my_reg[23][1]~q ;
wire \Mux30~7_combout ;
wire \Mux30~8_combout ;
wire \my_reg[3][1]~q ;
wire \my_reg[1][1]~feeder_combout ;
wire \my_reg[1][1]~q ;
wire \Mux30~14_combout ;
wire \my_reg[2][1]~q ;
wire \Mux30~15_combout ;
wire \my_reg[6][1]~q ;
wire \my_reg[7][1]~q ;
wire \my_reg[5][1]~q ;
wire \Decoder0~39_combout ;
wire \my_reg[4][1]~q ;
wire \Mux30~12_combout ;
wire \Mux30~13_combout ;
wire \Mux30~16_combout ;
wire \my_reg[9][1]~feeder_combout ;
wire \my_reg[9][1]~q ;
wire \my_reg[11][1]~q ;
wire \my_reg[10][1]~feeder_combout ;
wire \my_reg[10][1]~q ;
wire \Decoder0~33_combout ;
wire \my_reg[8][1]~q ;
wire \Mux30~10_combout ;
wire \Mux30~11_combout ;
wire \my_reg[15][1]~q ;
wire \my_reg[14][1]~q ;
wire \my_reg[13][1]~feeder_combout ;
wire \my_reg[13][1]~q ;
wire \Mux30~17_combout ;
wire \Mux30~18_combout ;
wire \my_reg[31][31]~q ;
wire \my_reg[27][31]~q ;
wire \my_reg[19][31]~feeder_combout ;
wire \Decoder0~29_combout ;
wire \my_reg[19][31]~q ;
wire \Mux0~7_combout ;
wire \Mux0~8_combout ;
wire \my_reg[25][31]~feeder_combout ;
wire \my_reg[25][31]~q ;
wire \my_reg[29][31]~q ;
wire \my_reg[21][31]~feeder_combout ;
wire \my_reg[21][31]~q ;
wire \my_reg[17][31]~feeder_combout ;
wire \Decoder0~14_combout ;
wire \my_reg[17][31]~q ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Decoder0~25_combout ;
wire \my_reg[28][31]~q ;
wire \my_reg[20][31]~q ;
wire \Mux0~5_combout ;
wire \my_reg[30][31]~q ;
wire \my_reg[18][31]~q ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \Mux0~6_combout ;
wire \Mux0~9_combout ;
wire \my_reg[9][31]~q ;
wire \my_reg[11][31]~q ;
wire \my_reg[8][31]~q ;
wire \Mux0~10_combout ;
wire \Mux0~11_combout ;
wire \my_reg[15][31]~q ;
wire \my_reg[13][31]~q ;
wire \my_reg[12][31]~q ;
wire \Mux0~17_combout ;
wire \Mux0~18_combout ;
wire \my_reg[2][31]~q ;
wire \my_reg[3][31]~q ;
wire \my_reg[1][31]~q ;
wire \Mux0~14_combout ;
wire \Mux0~15_combout ;
wire \my_reg[7][31]~q ;
wire \my_reg[4][31]~feeder_combout ;
wire \my_reg[4][31]~q ;
wire \Mux0~12_combout ;
wire \Mux0~13_combout ;
wire \Mux0~16_combout ;
wire \Mux0~19_combout ;
wire \my_reg[6][31]~feeder_combout ;
wire \my_reg[6][31]~q ;
wire \Mux32~0_combout ;
wire \Mux32~1_combout ;
wire \my_reg[14][31]~feeder_combout ;
wire \my_reg[14][31]~q ;
wire \Mux32~7_combout ;
wire \Mux32~8_combout ;
wire \Mux32~3_combout ;
wire \Mux32~4_combout ;
wire \Mux32~5_combout ;
wire \Mux32~6_combout ;
wire \my_reg[23][31]~feeder_combout ;
wire \my_reg[23][31]~q ;
wire \Mux32~17_combout ;
wire \Mux32~18_combout ;
wire \Mux32~10_combout ;
wire \Mux32~11_combout ;
wire \my_reg[24][31]~q ;
wire \my_reg[16][31]~q ;
wire \Mux32~14_combout ;
wire \Mux32~15_combout ;
wire \my_reg[26][31]~q ;
wire \Decoder0~18_combout ;
wire \my_reg[22][31]~q ;
wire \Mux32~12_combout ;
wire \Mux32~13_combout ;
wire \Mux32~16_combout ;
wire \my_reg[31][30]~q ;
wire \my_reg[19][30]~q ;
wire \Mux1~7_combout ;
wire \Mux1~8_combout ;
wire \my_reg[22][30]~q ;
wire \my_reg[18][30]~q ;
wire \Mux1~2_combout ;
wire \my_reg[30][30]~q ;
wire \Mux1~3_combout ;
wire \my_reg[24][30]~q ;
wire \my_reg[28][30]~q ;
wire \my_reg[20][30]~q ;
wire \my_reg[16][30]~q ;
wire \Mux1~4_combout ;
wire \Mux1~5_combout ;
wire \Mux1~6_combout ;
wire \my_reg[21][30]~feeder_combout ;
wire \my_reg[21][30]~q ;
wire \my_reg[29][30]~q ;
wire \my_reg[25][30]~feeder_combout ;
wire \my_reg[25][30]~q ;
wire \my_reg[17][30]~q ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux1~9_combout ;
wire \my_reg[9][30]~q ;
wire \my_reg[11][30]~q ;
wire \my_reg[8][30]~q ;
wire \Mux1~12_combout ;
wire \Mux1~13_combout ;
wire \my_reg[2][30]~feeder_combout ;
wire \my_reg[2][30]~q ;
wire \my_reg[1][30]~q ;
wire \my_reg[3][30]~q ;
wire \Mux1~14_combout ;
wire \Mux1~15_combout ;
wire \Mux1~16_combout ;
wire \my_reg[15][30]~q ;
wire \my_reg[13][30]~feeder_combout ;
wire \my_reg[13][30]~q ;
wire \my_reg[12][30]~q ;
wire \Mux1~17_combout ;
wire \Mux1~18_combout ;
wire \my_reg[6][30]~feeder_combout ;
wire \my_reg[6][30]~q ;
wire \my_reg[7][30]~q ;
wire \my_reg[5][30]~feeder_combout ;
wire \my_reg[5][30]~q ;
wire \Mux1~10_combout ;
wire \Mux1~11_combout ;
wire \Mux1~19_combout ;
wire \Mux33~0_combout ;
wire \Mux33~1_combout ;
wire \my_reg[4][30]~q ;
wire \Mux33~2_combout ;
wire \Mux33~3_combout ;
wire \Mux33~4_combout ;
wire \Mux33~5_combout ;
wire \Mux33~6_combout ;
wire \my_reg[14][30]~q ;
wire \Mux33~7_combout ;
wire \Mux33~8_combout ;
wire \Mux33~10_combout ;
wire \Mux33~11_combout ;
wire \my_reg[27][30]~q ;
wire \my_reg[23][30]~q ;
wire \Mux33~17_combout ;
wire \Mux33~18_combout ;
wire \Mux33~14_combout ;
wire \Mux33~15_combout ;
wire \my_reg[26][30]~q ;
wire \Mux33~12_combout ;
wire \Mux33~13_combout ;
wire \Mux33~16_combout ;
wire \my_reg[6][29]~q ;
wire \my_reg[7][29]~q ;
wire \my_reg[5][29]~q ;
wire \my_reg[4][29]~q ;
wire \Mux2~12_combout ;
wire \Mux2~13_combout ;
wire \my_reg[2][29]~q ;
wire \my_reg[3][29]~q ;
wire \Mux2~14_combout ;
wire \Mux2~15_combout ;
wire \Mux2~16_combout ;
wire \my_reg[10][29]~q ;
wire \my_reg[8][29]~q ;
wire \Mux2~10_combout ;
wire \my_reg[11][29]~q ;
wire \Mux2~11_combout ;
wire \my_reg[15][29]~q ;
wire \my_reg[13][29]~q ;
wire \my_reg[12][29]~q ;
wire \Mux2~17_combout ;
wire \Mux2~18_combout ;
wire \Mux2~19_combout ;
wire \my_reg[27][29]~q ;
wire \my_reg[31][29]~q ;
wire \my_reg[19][29]~q ;
wire \Mux2~7_combout ;
wire \Mux2~8_combout ;
wire \my_reg[25][29]~feeder_combout ;
wire \my_reg[25][29]~q ;
wire \my_reg[21][29]~feeder_combout ;
wire \my_reg[21][29]~q ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \my_reg[20][29]~q ;
wire \my_reg[28][29]~q ;
wire \my_reg[24][29]~feeder_combout ;
wire \my_reg[24][29]~q ;
wire \my_reg[16][29]~q ;
wire \Mux2~4_combout ;
wire \Mux2~5_combout ;
wire \my_reg[30][29]~q ;
wire \my_reg[26][29]~q ;
wire \Mux2~2_combout ;
wire \Mux2~3_combout ;
wire \Mux2~6_combout ;
wire \Mux2~9_combout ;
wire \Mux34~0_combout ;
wire \Mux34~1_combout ;
wire \my_reg[14][29]~q ;
wire \Mux34~7_combout ;
wire \Mux34~8_combout ;
wire \Mux34~2_combout ;
wire \my_reg[9][29]~q ;
wire \Mux34~3_combout ;
wire \my_reg[1][29]~feeder_combout ;
wire \my_reg[1][29]~q ;
wire \Mux34~4_combout ;
wire \Mux34~5_combout ;
wire \Mux34~6_combout ;
wire \Mux34~10_combout ;
wire \my_reg[29][29]~q ;
wire \Mux34~11_combout ;
wire \my_reg[18][29]~feeder_combout ;
wire \my_reg[18][29]~q ;
wire \my_reg[22][29]~q ;
wire \Mux34~12_combout ;
wire \Mux34~13_combout ;
wire \Mux34~14_combout ;
wire \Mux34~15_combout ;
wire \Mux34~16_combout ;
wire \my_reg[23][29]~feeder_combout ;
wire \my_reg[23][29]~q ;
wire \Mux34~17_combout ;
wire \Mux34~18_combout ;
wire \my_reg[2][28]~q ;
wire \my_reg[1][28]~q ;
wire \my_reg[3][28]~q ;
wire \Mux3~14_combout ;
wire \Mux3~15_combout ;
wire \my_reg[9][28]~q ;
wire \my_reg[11][28]~q ;
wire \my_reg[10][28]~q ;
wire \my_reg[8][28]~q ;
wire \Mux3~12_combout ;
wire \Mux3~13_combout ;
wire \Mux3~16_combout ;
wire \my_reg[15][28]~q ;
wire \my_reg[14][28]~q ;
wire \Mux3~18_combout ;
wire \my_reg[6][28]~q ;
wire \my_reg[7][28]~q ;
wire \my_reg[5][28]~q ;
wire \my_reg[4][28]~q ;
wire \Mux3~10_combout ;
wire \Mux3~11_combout ;
wire \Mux3~19_combout ;
wire \my_reg[19][28]~q ;
wire \Mux3~7_combout ;
wire \my_reg[31][28]~q ;
wire \Mux3~8_combout ;
wire \my_reg[26][28]~q ;
wire \my_reg[30][28]~q ;
wire \my_reg[18][28]~feeder_combout ;
wire \my_reg[18][28]~q ;
wire \my_reg[22][28]~q ;
wire \Mux3~2_combout ;
wire \Mux3~3_combout ;
wire \my_reg[24][28]~q ;
wire \my_reg[28][28]~q ;
wire \my_reg[20][28]~q ;
wire \my_reg[16][28]~q ;
wire \Mux3~4_combout ;
wire \Mux3~5_combout ;
wire \Mux3~6_combout ;
wire \my_reg[29][28]~q ;
wire \my_reg[17][28]~q ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Mux3~9_combout ;
wire \my_reg[13][28]~q ;
wire \Mux35~7_combout ;
wire \Mux35~8_combout ;
wire \Mux35~4_combout ;
wire \Mux35~5_combout ;
wire \Mux35~2_combout ;
wire \Mux35~3_combout ;
wire \Mux35~6_combout ;
wire \Mux35~0_combout ;
wire \Mux35~1_combout ;
wire \my_reg[25][28]~feeder_combout ;
wire \my_reg[25][28]~q ;
wire \Mux35~10_combout ;
wire \Mux35~11_combout ;
wire \my_reg[27][28]~q ;
wire \my_reg[23][28]~feeder_combout ;
wire \my_reg[23][28]~q ;
wire \Mux35~17_combout ;
wire \Mux35~18_combout ;
wire \Mux35~14_combout ;
wire \Mux35~15_combout ;
wire \Mux35~12_combout ;
wire \Mux35~13_combout ;
wire \Mux35~16_combout ;
wire \my_reg[25][27]~q ;
wire \my_reg[29][27]~q ;
wire \my_reg[17][27]~q ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;
wire \my_reg[22][27]~feeder_combout ;
wire \my_reg[22][27]~q ;
wire \my_reg[26][27]~feeder_combout ;
wire \my_reg[26][27]~q ;
wire \my_reg[18][27]~feeder_combout ;
wire \my_reg[18][27]~q ;
wire \Mux4~2_combout ;
wire \Mux4~3_combout ;
wire \my_reg[28][27]~feeder_combout ;
wire \my_reg[28][27]~q ;
wire \my_reg[16][27]~feeder_combout ;
wire \my_reg[16][27]~q ;
wire \Mux4~4_combout ;
wire \Mux4~5_combout ;
wire \Mux4~6_combout ;
wire \my_reg[27][27]~q ;
wire \my_reg[31][27]~q ;
wire \my_reg[19][27]~q ;
wire \Mux4~7_combout ;
wire \Mux4~8_combout ;
wire \Mux4~9_combout ;
wire \my_reg[15][27]~q ;
wire \my_reg[13][27]~feeder_combout ;
wire \my_reg[13][27]~q ;
wire \my_reg[12][27]~q ;
wire \Mux4~17_combout ;
wire \Mux4~18_combout ;
wire \my_reg[9][27]~feeder_combout ;
wire \my_reg[9][27]~q ;
wire \my_reg[10][27]~feeder_combout ;
wire \my_reg[10][27]~q ;
wire \Mux4~10_combout ;
wire \Mux4~11_combout ;
wire \my_reg[7][27]~feeder_combout ;
wire \my_reg[7][27]~q ;
wire \my_reg[6][27]~feeder_combout ;
wire \my_reg[6][27]~q ;
wire \my_reg[4][27]~feeder_combout ;
wire \my_reg[4][27]~q ;
wire \Mux4~12_combout ;
wire \Mux4~13_combout ;
wire \my_reg[2][27]~q ;
wire \my_reg[1][27]~q ;
wire \Mux4~14_combout ;
wire \Mux4~15_combout ;
wire \Mux4~16_combout ;
wire \Mux4~19_combout ;
wire \my_reg[14][27]~q ;
wire \Mux36~7_combout ;
wire \Mux36~8_combout ;
wire \my_reg[5][27]~feeder_combout ;
wire \my_reg[5][27]~q ;
wire \Mux36~0_combout ;
wire \Mux36~1_combout ;
wire \my_reg[11][27]~q ;
wire \my_reg[8][27]~q ;
wire \Mux36~2_combout ;
wire \Mux36~3_combout ;
wire \my_reg[3][27]~q ;
wire \Mux36~4_combout ;
wire \Mux36~5_combout ;
wire \Mux36~6_combout ;
wire \Mux36~10_combout ;
wire \my_reg[21][27]~feeder_combout ;
wire \my_reg[21][27]~q ;
wire \Mux36~11_combout ;
wire \my_reg[23][27]~q ;
wire \Mux36~17_combout ;
wire \Mux36~18_combout ;
wire \my_reg[24][27]~q ;
wire \my_reg[20][27]~q ;
wire \Mux36~14_combout ;
wire \Mux36~15_combout ;
wire \my_reg[30][27]~q ;
wire \Mux36~12_combout ;
wire \Mux36~13_combout ;
wire \Mux36~16_combout ;
wire \my_reg[31][26]~q ;
wire \my_reg[19][26]~q ;
wire \Mux5~7_combout ;
wire \Mux5~8_combout ;
wire \my_reg[21][26]~feeder_combout ;
wire \my_reg[21][26]~q ;
wire \my_reg[17][26]~q ;
wire \Mux5~0_combout ;
wire \my_reg[29][26]~feeder_combout ;
wire \my_reg[29][26]~q ;
wire \Mux5~1_combout ;
wire \my_reg[26][26]~q ;
wire \my_reg[30][26]~q ;
wire \my_reg[18][26]~feeder_combout ;
wire \my_reg[18][26]~q ;
wire \Mux5~2_combout ;
wire \Mux5~3_combout ;
wire \my_reg[24][26]~q ;
wire \my_reg[28][26]~q ;
wire \Mux5~5_combout ;
wire \Mux5~6_combout ;
wire \Mux5~9_combout ;
wire \my_reg[4][26]~q ;
wire \Mux5~10_combout ;
wire \my_reg[6][26]~feeder_combout ;
wire \my_reg[6][26]~q ;
wire \Mux5~11_combout ;
wire \my_reg[11][26]~q ;
wire \my_reg[10][26]~feeder_combout ;
wire \my_reg[10][26]~q ;
wire \my_reg[8][26]~q ;
wire \Mux5~12_combout ;
wire \Mux5~13_combout ;
wire \my_reg[3][26]~q ;
wire \my_reg[1][26]~q ;
wire \Mux5~14_combout ;
wire \Mux5~15_combout ;
wire \Mux5~16_combout ;
wire \my_reg[15][26]~feeder_combout ;
wire \my_reg[15][26]~q ;
wire \my_reg[13][26]~q ;
wire \my_reg[12][26]~q ;
wire \Mux5~17_combout ;
wire \Mux5~18_combout ;
wire \Mux5~19_combout ;
wire \my_reg[14][26]~q ;
wire \Mux37~7_combout ;
wire \Mux37~8_combout ;
wire \my_reg[9][26]~feeder_combout ;
wire \my_reg[9][26]~q ;
wire \Mux37~0_combout ;
wire \Mux37~1_combout ;
wire \Mux37~4_combout ;
wire \Mux37~5_combout ;
wire \my_reg[7][26]~q ;
wire \my_reg[5][26]~feeder_combout ;
wire \my_reg[5][26]~q ;
wire \Mux37~2_combout ;
wire \Mux37~3_combout ;
wire \Mux37~6_combout ;
wire \my_reg[27][26]~feeder_combout ;
wire \my_reg[27][26]~q ;
wire \Mux37~17_combout ;
wire \Mux37~18_combout ;
wire \my_reg[25][26]~feeder_combout ;
wire \my_reg[25][26]~q ;
wire \Mux37~10_combout ;
wire \Mux37~11_combout ;
wire \my_reg[20][26]~q ;
wire \my_reg[16][26]~q ;
wire \Mux37~14_combout ;
wire \Mux37~15_combout ;
wire \my_reg[22][26]~q ;
wire \Mux37~12_combout ;
wire \Mux37~13_combout ;
wire \Mux37~16_combout ;
wire \my_reg[9][25]~q ;
wire \my_reg[11][25]~q ;
wire \my_reg[10][25]~q ;
wire \my_reg[8][25]~q ;
wire \Mux6~10_combout ;
wire \Mux6~11_combout ;
wire \my_reg[14][25]~q ;
wire \my_reg[15][25]~q ;
wire \my_reg[13][25]~q ;
wire \my_reg[12][25]~q ;
wire \Mux6~17_combout ;
wire \Mux6~18_combout ;
wire \my_reg[6][25]~q ;
wire \my_reg[7][25]~q ;
wire \my_reg[4][25]~q ;
wire \my_reg[5][25]~q ;
wire \Mux6~12_combout ;
wire \Mux6~13_combout ;
wire \my_reg[2][25]~q ;
wire \Mux6~15_combout ;
wire \Mux6~16_combout ;
wire \Mux6~19_combout ;
wire \my_reg[29][25]~q ;
wire \my_reg[25][25]~q ;
wire \my_reg[17][25]~q ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \my_reg[20][25]~q ;
wire \my_reg[28][25]~q ;
wire \my_reg[24][25]~q ;
wire \my_reg[16][25]~q ;
wire \Mux6~4_combout ;
wire \Mux6~5_combout ;
wire \my_reg[30][25]~q ;
wire \my_reg[26][25]~q ;
wire \Mux6~2_combout ;
wire \Mux6~3_combout ;
wire \Mux6~6_combout ;
wire \my_reg[27][25]~q ;
wire \my_reg[31][25]~q ;
wire \my_reg[23][25]~q ;
wire \Mux6~7_combout ;
wire \Mux6~8_combout ;
wire \Mux6~9_combout ;
wire \my_reg[3][25]~q ;
wire \Mux38~4_combout ;
wire \Mux38~5_combout ;
wire \Mux38~2_combout ;
wire \Mux38~3_combout ;
wire \Mux38~6_combout ;
wire \Mux38~7_combout ;
wire \Mux38~8_combout ;
wire \Mux38~0_combout ;
wire \Mux38~1_combout ;
wire \my_reg[21][25]~feeder_combout ;
wire \my_reg[21][25]~q ;
wire \Mux38~10_combout ;
wire \Mux38~11_combout ;
wire \my_reg[19][25]~feeder_combout ;
wire \my_reg[19][25]~q ;
wire \Mux38~17_combout ;
wire \Mux38~18_combout ;
wire \Mux38~14_combout ;
wire \Mux38~15_combout ;
wire \my_reg[18][25]~feeder_combout ;
wire \my_reg[18][25]~q ;
wire \my_reg[22][25]~q ;
wire \Mux38~12_combout ;
wire \Mux38~13_combout ;
wire \Mux38~16_combout ;
wire \my_reg[21][24]~feeder_combout ;
wire \my_reg[21][24]~q ;
wire \my_reg[29][24]~q ;
wire \my_reg[25][24]~feeder_combout ;
wire \my_reg[25][24]~q ;
wire \my_reg[17][24]~q ;
wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \my_reg[23][24]~q ;
wire \my_reg[31][24]~q ;
wire \my_reg[19][24]~q ;
wire \Mux7~7_combout ;
wire \Mux7~8_combout ;
wire \my_reg[24][24]~q ;
wire \my_reg[28][24]~q ;
wire \my_reg[16][24]~q ;
wire \Mux7~4_combout ;
wire \Mux7~5_combout ;
wire \my_reg[30][24]~q ;
wire \my_reg[18][24]~q ;
wire \Mux7~2_combout ;
wire \Mux7~3_combout ;
wire \Mux7~6_combout ;
wire \my_reg[7][24]~q ;
wire \my_reg[6][24]~q ;
wire \my_reg[4][24]~q ;
wire \my_reg[5][24]~q ;
wire \Mux7~10_combout ;
wire \Mux7~11_combout ;
wire \my_reg[15][24]~q ;
wire \my_reg[14][24]~feeder_combout ;
wire \my_reg[14][24]~q ;
wire \my_reg[12][24]~feeder_combout ;
wire \my_reg[12][24]~q ;
wire \my_reg[13][24]~q ;
wire \Mux7~17_combout ;
wire \Mux7~18_combout ;
wire \my_reg[9][24]~q ;
wire \my_reg[11][24]~q ;
wire \my_reg[10][24]~q ;
wire \my_reg[8][24]~q ;
wire \Mux7~12_combout ;
wire \Mux7~13_combout ;
wire \my_reg[2][24]~q ;
wire \my_reg[1][24]~q ;
wire \Mux7~14_combout ;
wire \Mux7~15_combout ;
wire \Mux7~16_combout ;
wire \my_reg[3][24]~q ;
wire \Mux39~4_combout ;
wire \Mux39~5_combout ;
wire \Mux39~2_combout ;
wire \Mux39~3_combout ;
wire \Mux39~6_combout ;
wire \Mux39~7_combout ;
wire \Mux39~8_combout ;
wire \Mux39~0_combout ;
wire \Mux39~1_combout ;
wire \Mux39~10_combout ;
wire \Mux39~11_combout ;
wire \my_reg[27][24]~q ;
wire \Mux39~17_combout ;
wire \Mux39~18_combout ;
wire \Mux39~14_combout ;
wire \my_reg[20][24]~q ;
wire \Mux39~15_combout ;
wire \my_reg[22][24]~q ;
wire \my_reg[26][24]~q ;
wire \Mux39~12_combout ;
wire \Mux39~13_combout ;
wire \Mux39~16_combout ;
wire \my_reg[11][23]~q ;
wire \my_reg[9][23]~feeder_combout ;
wire \my_reg[9][23]~q ;
wire \Mux8~11_combout ;
wire \my_reg[14][23]~q ;
wire \my_reg[15][23]~q ;
wire \my_reg[12][23]~feeder_combout ;
wire \my_reg[12][23]~q ;
wire \Mux8~17_combout ;
wire \Mux8~18_combout ;
wire \my_reg[6][23]~q ;
wire \my_reg[7][23]~q ;
wire \my_reg[4][23]~feeder_combout ;
wire \my_reg[4][23]~q ;
wire \Mux8~12_combout ;
wire \Mux8~13_combout ;
wire \my_reg[3][23]~q ;
wire \my_reg[1][23]~q ;
wire \Mux8~14_combout ;
wire \my_reg[2][23]~q ;
wire \Mux8~15_combout ;
wire \Mux8~16_combout ;
wire \Mux8~19_combout ;
wire \my_reg[27][23]~q ;
wire \my_reg[31][23]~q ;
wire \my_reg[23][23]~q ;
wire \my_reg[19][23]~q ;
wire \Mux8~7_combout ;
wire \Mux8~8_combout ;
wire \my_reg[25][23]~feeder_combout ;
wire \my_reg[25][23]~q ;
wire \my_reg[29][23]~q ;
wire \my_reg[17][23]~q ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \my_reg[28][23]~q ;
wire \my_reg[16][23]~q ;
wire \Mux8~4_combout ;
wire \Mux8~5_combout ;
wire \my_reg[22][23]~q ;
wire \my_reg[30][23]~q ;
wire \my_reg[26][23]~q ;
wire \my_reg[18][23]~q ;
wire \Mux8~2_combout ;
wire \Mux8~3_combout ;
wire \Mux8~6_combout ;
wire \Mux8~9_combout ;
wire \my_reg[5][23]~q ;
wire \Mux40~0_combout ;
wire \Mux40~1_combout ;
wire \my_reg[10][23]~feeder_combout ;
wire \my_reg[10][23]~q ;
wire \my_reg[8][23]~q ;
wire \Mux40~2_combout ;
wire \Mux40~3_combout ;
wire \Mux40~4_combout ;
wire \Mux40~5_combout ;
wire \Mux40~6_combout ;
wire \Mux40~7_combout ;
wire \Mux40~8_combout ;
wire \Mux40~17_combout ;
wire \Mux40~18_combout ;
wire \Mux40~10_combout ;
wire \my_reg[21][23]~q ;
wire \Mux40~11_combout ;
wire \my_reg[24][23]~q ;
wire \my_reg[20][23]~q ;
wire \Mux40~14_combout ;
wire \Mux40~15_combout ;
wire \Mux40~12_combout ;
wire \Mux40~13_combout ;
wire \Mux40~16_combout ;
wire \my_reg[15][22]~feeder_combout ;
wire \my_reg[15][22]~q ;
wire \my_reg[13][22]~q ;
wire \my_reg[12][22]~q ;
wire \Mux9~17_combout ;
wire \Mux9~18_combout ;
wire \my_reg[6][22]~q ;
wire \my_reg[7][22]~q ;
wire \my_reg[4][22]~q ;
wire \Mux9~10_combout ;
wire \Mux9~11_combout ;
wire \my_reg[2][22]~q ;
wire \my_reg[1][22]~q ;
wire \Mux9~14_combout ;
wire \Mux9~15_combout ;
wire \my_reg[9][22]~q ;
wire \my_reg[11][22]~q ;
wire \my_reg[10][22]~feeder_combout ;
wire \my_reg[10][22]~q ;
wire \my_reg[8][22]~q ;
wire \Mux9~12_combout ;
wire \Mux9~13_combout ;
wire \Mux9~16_combout ;
wire \Mux9~19_combout ;
wire \my_reg[23][22]~q ;
wire \my_reg[31][22]~q ;
wire \my_reg[27][22]~q ;
wire \my_reg[19][22]~q ;
wire \Mux9~7_combout ;
wire \Mux9~8_combout ;
wire \my_reg[21][22]~q ;
wire \my_reg[29][22]~q ;
wire \my_reg[17][22]~q ;
wire \Mux9~0_combout ;
wire \Mux9~1_combout ;
wire \my_reg[30][22]~q ;
wire \my_reg[18][22]~q ;
wire \Mux9~2_combout ;
wire \Mux9~3_combout ;
wire \my_reg[28][22]~q ;
wire \my_reg[16][22]~q ;
wire \my_reg[20][22]~q ;
wire \Mux9~4_combout ;
wire \Mux9~5_combout ;
wire \Mux9~6_combout ;
wire \Mux9~9_combout ;
wire \Mux41~0_combout ;
wire \Mux41~1_combout ;
wire \Mux41~5_combout ;
wire \Mux41~3_combout ;
wire \Mux41~6_combout ;
wire \Mux41~7_combout ;
wire \my_reg[14][22]~q ;
wire \Mux41~8_combout ;
wire \Mux41~17_combout ;
wire \Mux41~18_combout ;
wire \my_reg[25][22]~feeder_combout ;
wire \my_reg[25][22]~q ;
wire \Mux41~10_combout ;
wire \Mux41~11_combout ;
wire \my_reg[24][22]~q ;
wire \Mux41~14_combout ;
wire \Mux41~15_combout ;
wire \my_reg[22][22]~q ;
wire \my_reg[26][22]~q ;
wire \Mux41~12_combout ;
wire \Mux41~13_combout ;
wire \Mux41~16_combout ;
wire \my_reg[2][21]~q ;
wire \Mux10~15_combout ;
wire \my_reg[6][21]~q ;
wire \my_reg[7][21]~q ;
wire \my_reg[4][21]~feeder_combout ;
wire \my_reg[4][21]~q ;
wire \Mux10~12_combout ;
wire \Mux10~13_combout ;
wire \Mux10~16_combout ;
wire \my_reg[15][21]~q ;
wire \my_reg[14][21]~q ;
wire \Mux10~18_combout ;
wire \my_reg[9][21]~q ;
wire \my_reg[11][21]~q ;
wire \my_reg[10][21]~q ;
wire \my_reg[8][21]~feeder_combout ;
wire \my_reg[8][21]~q ;
wire \Mux10~10_combout ;
wire \Mux10~11_combout ;
wire \Mux10~19_combout ;
wire \my_reg[27][21]~q ;
wire \my_reg[31][21]~q ;
wire \my_reg[19][21]~q ;
wire \Mux10~7_combout ;
wire \Mux10~8_combout ;
wire \my_reg[25][21]~q ;
wire \my_reg[29][21]~q ;
wire \my_reg[21][21]~q ;
wire \my_reg[17][21]~q ;
wire \Mux10~0_combout ;
wire \Mux10~1_combout ;
wire \my_reg[30][21]~feeder_combout ;
wire \my_reg[30][21]~q ;
wire \my_reg[18][21]~feeder_combout ;
wire \my_reg[18][21]~q ;
wire \my_reg[26][21]~q ;
wire \Mux10~2_combout ;
wire \Mux10~3_combout ;
wire \my_reg[20][21]~q ;
wire \my_reg[28][21]~q ;
wire \my_reg[24][21]~feeder_combout ;
wire \my_reg[24][21]~q ;
wire \my_reg[16][21]~feeder_combout ;
wire \my_reg[16][21]~q ;
wire \Mux10~4_combout ;
wire \Mux10~5_combout ;
wire \Mux10~6_combout ;
wire \Mux10~9_combout ;
wire \my_reg[3][21]~q ;
wire \Mux42~4_combout ;
wire \Mux42~5_combout ;
wire \Mux42~3_combout ;
wire \Mux42~6_combout ;
wire \my_reg[5][21]~q ;
wire \Mux42~0_combout ;
wire \Mux42~1_combout ;
wire \my_reg[13][21]~q ;
wire \Mux42~7_combout ;
wire \Mux42~8_combout ;
wire \Mux42~10_combout ;
wire \Mux42~11_combout ;
wire \Mux42~14_combout ;
wire \Mux42~15_combout ;
wire \my_reg[22][21]~q ;
wire \Mux42~12_combout ;
wire \Mux42~13_combout ;
wire \Mux42~16_combout ;
wire \my_reg[23][21]~q ;
wire \Mux42~17_combout ;
wire \Mux42~18_combout ;
wire \my_reg[2][20]~q ;
wire \my_reg[1][20]~q ;
wire \Mux11~14_combout ;
wire \Mux11~15_combout ;
wire \Mux11~16_combout ;
wire \my_reg[6][20]~q ;
wire \my_reg[5][20]~q ;
wire \my_reg[4][20]~q ;
wire \Mux11~10_combout ;
wire \Mux11~11_combout ;
wire \my_reg[14][20]~q ;
wire \my_reg[15][20]~q ;
wire \my_reg[13][20]~q ;
wire \my_reg[12][20]~q ;
wire \Mux11~17_combout ;
wire \Mux11~18_combout ;
wire \Mux11~19_combout ;
wire \my_reg[23][20]~q ;
wire \my_reg[31][20]~q ;
wire \my_reg[27][20]~q ;
wire \my_reg[19][20]~q ;
wire \Mux11~7_combout ;
wire \Mux11~8_combout ;
wire \my_reg[21][20]~q ;
wire \my_reg[17][20]~q ;
wire \my_reg[25][20]~feeder_combout ;
wire \my_reg[25][20]~q ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \my_reg[30][20]~q ;
wire \my_reg[18][20]~q ;
wire \Mux11~2_combout ;
wire \Mux11~3_combout ;
wire \my_reg[28][20]~q ;
wire \my_reg[20][20]~q ;
wire \Mux11~4_combout ;
wire \Mux11~5_combout ;
wire \Mux11~6_combout ;
wire \Mux11~9_combout ;
wire \my_reg[8][20]~q ;
wire \my_reg[10][20]~q ;
wire \Mux43~0_combout ;
wire \my_reg[11][20]~q ;
wire \my_reg[9][20]~q ;
wire \Mux43~1_combout ;
wire \my_reg[7][20]~feeder_combout ;
wire \my_reg[7][20]~q ;
wire \Mux43~2_combout ;
wire \Mux43~3_combout ;
wire \my_reg[3][20]~q ;
wire \Mux43~4_combout ;
wire \Mux43~5_combout ;
wire \Mux43~6_combout ;
wire \Mux43~7_combout ;
wire \Mux43~8_combout ;
wire \Mux43~17_combout ;
wire \Mux43~18_combout ;
wire \Mux43~10_combout ;
wire \my_reg[29][20]~feeder_combout ;
wire \my_reg[29][20]~q ;
wire \Mux43~11_combout ;
wire \my_reg[16][20]~q ;
wire \my_reg[24][20]~q ;
wire \Mux43~14_combout ;
wire \Mux43~15_combout ;
wire \my_reg[22][20]~feeder_combout ;
wire \my_reg[22][20]~q ;
wire \my_reg[26][20]~q ;
wire \Mux43~12_combout ;
wire \Mux43~13_combout ;
wire \Mux43~16_combout ;
wire \my_reg[19][19]~q ;
wire \Mux12~7_combout ;
wire \my_reg[31][19]~q ;
wire \Mux12~8_combout ;
wire \my_reg[16][19]~q ;
wire \Mux12~4_combout ;
wire \my_reg[28][19]~q ;
wire \Mux12~5_combout ;
wire \my_reg[22][19]~q ;
wire \my_reg[30][19]~q ;
wire \my_reg[26][19]~q ;
wire \my_reg[18][19]~feeder_combout ;
wire \my_reg[18][19]~q ;
wire \Mux12~2_combout ;
wire \Mux12~3_combout ;
wire \Mux12~6_combout ;
wire \my_reg[25][19]~feeder_combout ;
wire \my_reg[25][19]~q ;
wire \my_reg[29][19]~q ;
wire \my_reg[17][19]~feeder_combout ;
wire \my_reg[17][19]~q ;
wire \Mux12~0_combout ;
wire \Mux12~1_combout ;
wire \Mux12~9_combout ;
wire \my_reg[15][19]~q ;
wire \my_reg[13][19]~q ;
wire \my_reg[12][19]~q ;
wire \Mux12~17_combout ;
wire \Mux12~18_combout ;
wire \my_reg[9][19]~q ;
wire \my_reg[11][19]~q ;
wire \my_reg[8][19]~q ;
wire \Mux12~10_combout ;
wire \Mux12~11_combout ;
wire \my_reg[7][19]~q ;
wire \my_reg[5][19]~q ;
wire \my_reg[4][19]~q ;
wire \Mux12~12_combout ;
wire \Mux12~13_combout ;
wire \my_reg[2][19]~q ;
wire \my_reg[1][19]~q ;
wire \Mux12~14_combout ;
wire \Mux12~15_combout ;
wire \Mux12~16_combout ;
wire \Mux12~19_combout ;
wire \my_reg[10][19]~q ;
wire \Mux44~2_combout ;
wire \Mux44~3_combout ;
wire \my_reg[3][19]~feeder_combout ;
wire \my_reg[3][19]~q ;
wire \Mux44~4_combout ;
wire \Mux44~5_combout ;
wire \Mux44~6_combout ;
wire \my_reg[14][19]~feeder_combout ;
wire \my_reg[14][19]~q ;
wire \Mux44~7_combout ;
wire \Mux44~8_combout ;
wire \Mux44~0_combout ;
wire \my_reg[6][19]~q ;
wire \Mux44~1_combout ;
wire \my_reg[21][19]~q ;
wire \Mux44~10_combout ;
wire \Mux44~11_combout ;
wire \Mux44~17_combout ;
wire \my_reg[23][19]~feeder_combout ;
wire \my_reg[23][19]~q ;
wire \Mux44~18_combout ;
wire \my_reg[24][19]~q ;
wire \my_reg[20][19]~q ;
wire \Mux44~14_combout ;
wire \Mux44~15_combout ;
wire \Mux44~12_combout ;
wire \Mux44~13_combout ;
wire \Mux44~16_combout ;
wire \my_reg[15][18]~q ;
wire \my_reg[14][18]~q ;
wire \my_reg[12][18]~q ;
wire \Mux13~17_combout ;
wire \Mux13~18_combout ;
wire \my_reg[4][18]~q ;
wire \Mux13~10_combout ;
wire \my_reg[7][18]~q ;
wire \Mux13~11_combout ;
wire \my_reg[2][18]~q ;
wire \my_reg[1][18]~q ;
wire \Mux13~14_combout ;
wire \Mux13~15_combout ;
wire \my_reg[9][18]~q ;
wire \my_reg[11][18]~q ;
wire \my_reg[8][18]~q ;
wire \Mux13~12_combout ;
wire \Mux13~13_combout ;
wire \Mux13~16_combout ;
wire \Mux13~19_combout ;
wire \my_reg[27][18]~q ;
wire \my_reg[19][18]~q ;
wire \Mux13~7_combout ;
wire \my_reg[31][18]~q ;
wire \Mux13~8_combout ;
wire \my_reg[30][18]~feeder_combout ;
wire \my_reg[30][18]~q ;
wire \my_reg[18][18]~q ;
wire \Mux13~2_combout ;
wire \Mux13~3_combout ;
wire \my_reg[16][18]~q ;
wire \Mux13~4_combout ;
wire \my_reg[28][18]~q ;
wire \Mux13~5_combout ;
wire \Mux13~6_combout ;
wire \my_reg[21][18]~feeder_combout ;
wire \my_reg[21][18]~q ;
wire \my_reg[29][18]~q ;
wire \my_reg[25][18]~feeder_combout ;
wire \my_reg[25][18]~q ;
wire \my_reg[17][18]~feeder_combout ;
wire \my_reg[17][18]~q ;
wire \Mux13~0_combout ;
wire \Mux13~1_combout ;
wire \Mux13~9_combout ;
wire \my_reg[13][18]~feeder_combout ;
wire \my_reg[13][18]~q ;
wire \Mux45~7_combout ;
wire \Mux45~8_combout ;
wire \my_reg[10][18]~q ;
wire \Mux45~0_combout ;
wire \Mux45~1_combout ;
wire \my_reg[3][18]~q ;
wire \Mux45~4_combout ;
wire \Mux45~5_combout ;
wire \my_reg[6][18]~q ;
wire \Mux45~3_combout ;
wire \Mux45~6_combout ;
wire \my_reg[23][18]~q ;
wire \Mux45~17_combout ;
wire \Mux45~18_combout ;
wire \my_reg[20][18]~q ;
wire \my_reg[24][18]~q ;
wire \Mux45~14_combout ;
wire \Mux45~15_combout ;
wire \my_reg[22][18]~feeder_combout ;
wire \my_reg[22][18]~q ;
wire \my_reg[26][18]~q ;
wire \Mux45~12_combout ;
wire \Mux45~13_combout ;
wire \Mux45~16_combout ;
wire \Mux45~10_combout ;
wire \Mux45~11_combout ;
wire \my_reg[6][17]~q ;
wire \my_reg[7][17]~q ;
wire \my_reg[5][17]~q ;
wire \Mux14~12_combout ;
wire \Mux14~13_combout ;
wire \my_reg[2][17]~q ;
wire \my_reg[1][17]~q ;
wire \Mux14~14_combout ;
wire \Mux14~15_combout ;
wire \Mux14~16_combout ;
wire \my_reg[15][17]~feeder_combout ;
wire \my_reg[15][17]~q ;
wire \my_reg[14][17]~q ;
wire \my_reg[12][17]~q ;
wire \Mux14~17_combout ;
wire \Mux14~18_combout ;
wire \my_reg[9][17]~feeder_combout ;
wire \my_reg[9][17]~q ;
wire \my_reg[10][17]~q ;
wire \Mux14~10_combout ;
wire \Mux14~11_combout ;
wire \Mux14~19_combout ;
wire \my_reg[27][17]~q ;
wire \my_reg[31][17]~q ;
wire \my_reg[23][17]~q ;
wire \my_reg[19][17]~q ;
wire \Mux14~7_combout ;
wire \Mux14~8_combout ;
wire \my_reg[25][17]~feeder_combout ;
wire \my_reg[25][17]~q ;
wire \my_reg[29][17]~q ;
wire \my_reg[17][17]~q ;
wire \my_reg[21][17]~feeder_combout ;
wire \my_reg[21][17]~q ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \my_reg[28][17]~q ;
wire \my_reg[16][17]~q ;
wire \Mux14~4_combout ;
wire \Mux14~5_combout ;
wire \my_reg[22][17]~q ;
wire \my_reg[30][17]~q ;
wire \my_reg[18][17]~feeder_combout ;
wire \my_reg[18][17]~q ;
wire \Mux14~2_combout ;
wire \Mux14~3_combout ;
wire \Mux14~6_combout ;
wire \Mux14~9_combout ;
wire \my_reg[4][17]~feeder_combout ;
wire \my_reg[4][17]~q ;
wire \Mux46~0_combout ;
wire \Mux46~1_combout ;
wire \my_reg[13][17]~feeder_combout ;
wire \my_reg[13][17]~q ;
wire \Mux46~7_combout ;
wire \Mux46~8_combout ;
wire \my_reg[3][17]~q ;
wire \Mux46~4_combout ;
wire \Mux46~5_combout ;
wire \my_reg[8][17]~q ;
wire \Mux46~2_combout ;
wire \my_reg[11][17]~q ;
wire \Mux46~3_combout ;
wire \Mux46~6_combout ;
wire \Mux46~10_combout ;
wire \Mux46~11_combout ;
wire \Mux46~17_combout ;
wire \Mux46~18_combout ;
wire \my_reg[24][17]~feeder_combout ;
wire \my_reg[24][17]~q ;
wire \Mux46~14_combout ;
wire \Mux46~15_combout ;
wire \my_reg[26][17]~q ;
wire \Mux46~12_combout ;
wire \Mux46~13_combout ;
wire \Mux46~16_combout ;
wire \my_reg[2][16]~q ;
wire \my_reg[1][16]~q ;
wire \my_reg[3][16]~q ;
wire \Mux15~14_combout ;
wire \Mux15~15_combout ;
wire \my_reg[9][16]~q ;
wire \my_reg[11][16]~q ;
wire \my_reg[10][16]~q ;
wire \my_reg[8][16]~q ;
wire \Mux15~12_combout ;
wire \Mux15~13_combout ;
wire \Mux15~16_combout ;
wire \my_reg[14][16]~q ;
wire \my_reg[15][16]~q ;
wire \my_reg[12][16]~q ;
wire \Mux15~17_combout ;
wire \Mux15~18_combout ;
wire \my_reg[7][16]~q ;
wire \my_reg[6][16]~q ;
wire \my_reg[4][16]~q ;
wire \my_reg[5][16]~q ;
wire \Mux15~10_combout ;
wire \Mux15~11_combout ;
wire \Mux15~19_combout ;
wire \my_reg[23][16]~feeder_combout ;
wire \my_reg[23][16]~q ;
wire \my_reg[31][16]~q ;
wire \my_reg[27][16]~feeder_combout ;
wire \my_reg[27][16]~q ;
wire \my_reg[19][16]~q ;
wire \Mux15~7_combout ;
wire \Mux15~8_combout ;
wire \my_reg[29][16]~q ;
wire \my_reg[25][16]~feeder_combout ;
wire \my_reg[25][16]~q ;
wire \my_reg[17][16]~q ;
wire \Mux15~0_combout ;
wire \Mux15~1_combout ;
wire \my_reg[24][16]~feeder_combout ;
wire \my_reg[24][16]~q ;
wire \my_reg[28][16]~q ;
wire \my_reg[16][16]~feeder_combout ;
wire \my_reg[16][16]~q ;
wire \Mux15~4_combout ;
wire \Mux15~5_combout ;
wire \Mux15~6_combout ;
wire \Mux15~9_combout ;
wire \Mux47~0_combout ;
wire \Mux47~1_combout ;
wire \my_reg[13][16]~q ;
wire \Mux47~7_combout ;
wire \Mux47~8_combout ;
wire \Mux47~2_combout ;
wire \Mux47~3_combout ;
wire \Mux47~4_combout ;
wire \Mux47~5_combout ;
wire \Mux47~6_combout ;
wire \my_reg[21][16]~q ;
wire \Mux47~10_combout ;
wire \Mux47~11_combout ;
wire \my_reg[22][16]~q ;
wire \my_reg[18][16]~q ;
wire \my_reg[26][16]~q ;
wire \Mux47~12_combout ;
wire \Mux47~13_combout ;
wire \my_reg[20][16]~q ;
wire \Mux47~14_combout ;
wire \Mux47~15_combout ;
wire \Mux47~16_combout ;
wire \Mux47~17_combout ;
wire \Mux47~18_combout ;
wire \my_reg[19][15]~q ;
wire \Mux16~7_combout ;
wire \my_reg[31][15]~q ;
wire \Mux16~8_combout ;
wire \my_reg[22][15]~q ;
wire \my_reg[30][15]~feeder_combout ;
wire \my_reg[30][15]~q ;
wire \my_reg[18][15]~feeder_combout ;
wire \my_reg[18][15]~q ;
wire \Mux16~2_combout ;
wire \Mux16~3_combout ;
wire \my_reg[28][15]~q ;
wire \my_reg[16][15]~q ;
wire \Mux16~4_combout ;
wire \Mux16~5_combout ;
wire \Mux16~6_combout ;
wire \my_reg[29][15]~feeder_combout ;
wire \my_reg[29][15]~q ;
wire \my_reg[17][15]~q ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \Mux16~9_combout ;
wire \my_reg[15][15]~feeder_combout ;
wire \my_reg[15][15]~q ;
wire \my_reg[12][15]~feeder_combout ;
wire \my_reg[12][15]~q ;
wire \my_reg[13][15]~q ;
wire \Mux16~17_combout ;
wire \Mux16~18_combout ;
wire \my_reg[9][15]~feeder_combout ;
wire \my_reg[9][15]~q ;
wire \my_reg[10][15]~q ;
wire \Mux16~10_combout ;
wire \my_reg[11][15]~q ;
wire \Mux16~11_combout ;
wire \my_reg[3][15]~q ;
wire \Mux16~14_combout ;
wire \Mux16~15_combout ;
wire \my_reg[7][15]~q ;
wire \my_reg[4][15]~q ;
wire \Mux16~12_combout ;
wire \Mux16~13_combout ;
wire \Mux16~16_combout ;
wire \Mux16~19_combout ;
wire \my_reg[5][15]~q ;
wire \Mux48~0_combout ;
wire \my_reg[6][15]~q ;
wire \Mux48~1_combout ;
wire \my_reg[14][15]~feeder_combout ;
wire \my_reg[14][15]~q ;
wire \Mux48~7_combout ;
wire \Mux48~8_combout ;
wire \my_reg[8][15]~q ;
wire \Mux48~2_combout ;
wire \Mux48~3_combout ;
wire \my_reg[2][15]~q ;
wire \my_reg[1][15]~q ;
wire \Mux48~4_combout ;
wire \Mux48~5_combout ;
wire \Mux48~6_combout ;
wire \my_reg[23][15]~feeder_combout ;
wire \my_reg[23][15]~q ;
wire \Mux48~17_combout ;
wire \Mux48~18_combout ;
wire \my_reg[24][15]~feeder_combout ;
wire \my_reg[24][15]~q ;
wire \Mux48~15_combout ;
wire \my_reg[26][15]~q ;
wire \Mux48~12_combout ;
wire \Mux48~13_combout ;
wire \Mux48~16_combout ;
wire \my_reg[21][15]~feeder_combout ;
wire \my_reg[21][15]~q ;
wire \my_reg[25][15]~feeder_combout ;
wire \my_reg[25][15]~q ;
wire \Mux48~10_combout ;
wire \Mux48~11_combout ;
wire \my_reg[14][14]~feeder_combout ;
wire \my_reg[14][14]~q ;
wire \my_reg[12][14]~q ;
wire \my_reg[13][14]~q ;
wire \Mux17~17_combout ;
wire \Mux17~18_combout ;
wire \my_reg[7][14]~feeder_combout ;
wire \my_reg[7][14]~q ;
wire \my_reg[4][14]~q ;
wire \Mux17~10_combout ;
wire \Mux17~11_combout ;
wire \my_reg[2][14]~q ;
wire \my_reg[1][14]~q ;
wire \my_reg[3][14]~q ;
wire \Mux17~14_combout ;
wire \Mux17~15_combout ;
wire \my_reg[9][14]~q ;
wire \my_reg[11][14]~q ;
wire \my_reg[8][14]~q ;
wire \Mux17~12_combout ;
wire \Mux17~13_combout ;
wire \Mux17~16_combout ;
wire \Mux17~19_combout ;
wire \my_reg[21][14]~q ;
wire \my_reg[29][14]~q ;
wire \Mux17~1_combout ;
wire \my_reg[31][14]~feeder_combout ;
wire \my_reg[31][14]~q ;
wire \my_reg[27][14]~q ;
wire \Mux17~7_combout ;
wire \Mux17~8_combout ;
wire \my_reg[28][14]~q ;
wire \my_reg[16][14]~q ;
wire \Mux17~4_combout ;
wire \Mux17~5_combout ;
wire \my_reg[26][14]~q ;
wire \my_reg[30][14]~feeder_combout ;
wire \my_reg[30][14]~q ;
wire \my_reg[18][14]~q ;
wire \Mux17~2_combout ;
wire \Mux17~3_combout ;
wire \Mux17~6_combout ;
wire \Mux17~9_combout ;
wire \my_reg[15][14]~feeder_combout ;
wire \my_reg[15][14]~q ;
wire \Mux49~7_combout ;
wire \Mux49~8_combout ;
wire \my_reg[10][14]~q ;
wire \Mux49~0_combout ;
wire \Mux49~1_combout ;
wire \my_reg[6][14]~feeder_combout ;
wire \my_reg[6][14]~q ;
wire \Mux49~2_combout ;
wire \Mux49~3_combout ;
wire \Mux49~4_combout ;
wire \Mux49~5_combout ;
wire \Mux49~6_combout ;
wire \my_reg[25][14]~feeder_combout ;
wire \my_reg[25][14]~q ;
wire \Mux49~10_combout ;
wire \Mux49~11_combout ;
wire \my_reg[20][14]~q ;
wire \Mux49~15_combout ;
wire \Mux49~12_combout ;
wire \my_reg[22][14]~q ;
wire \Mux49~13_combout ;
wire \Mux49~16_combout ;
wire \my_reg[19][14]~feeder_combout ;
wire \my_reg[19][14]~q ;
wire \my_reg[23][14]~q ;
wire \Mux49~17_combout ;
wire \Mux49~18_combout ;
wire \my_reg[9][13]~feeder_combout ;
wire \my_reg[9][13]~q ;
wire \my_reg[8][13]~q ;
wire \Mux18~10_combout ;
wire \Mux18~11_combout ;
wire \my_reg[2][13]~q ;
wire \Mux18~15_combout ;
wire \my_reg[6][13]~q ;
wire \my_reg[7][13]~q ;
wire \my_reg[4][13]~q ;
wire \Mux18~12_combout ;
wire \Mux18~13_combout ;
wire \Mux18~16_combout ;
wire \my_reg[14][13]~q ;
wire \my_reg[13][13]~feeder_combout ;
wire \my_reg[13][13]~q ;
wire \Mux18~17_combout ;
wire \Mux18~18_combout ;
wire \Mux18~19_combout ;
wire \my_reg[16][13]~q ;
wire \Mux18~4_combout ;
wire \my_reg[20][13]~q ;
wire \Mux18~5_combout ;
wire \Mux18~6_combout ;
wire \my_reg[29][13]~q ;
wire \my_reg[17][13]~feeder_combout ;
wire \my_reg[17][13]~q ;
wire \Mux18~0_combout ;
wire \Mux18~1_combout ;
wire \my_reg[27][13]~q ;
wire \my_reg[31][13]~q ;
wire \my_reg[19][13]~feeder_combout ;
wire \my_reg[19][13]~q ;
wire \Mux18~7_combout ;
wire \Mux18~8_combout ;
wire \Mux18~9_combout ;
wire \my_reg[15][13]~q ;
wire \Mux50~7_combout ;
wire \Mux50~8_combout ;
wire \my_reg[3][13]~q ;
wire \Mux50~4_combout ;
wire \Mux50~5_combout ;
wire \my_reg[11][13]~q ;
wire \my_reg[10][13]~feeder_combout ;
wire \my_reg[10][13]~q ;
wire \Mux50~2_combout ;
wire \Mux50~3_combout ;
wire \Mux50~6_combout ;
wire \my_reg[5][13]~q ;
wire \Mux50~0_combout ;
wire \Mux50~1_combout ;
wire \my_reg[21][13]~feeder_combout ;
wire \my_reg[21][13]~q ;
wire \my_reg[25][13]~q ;
wire \Mux50~10_combout ;
wire \Mux50~11_combout ;
wire \my_reg[23][13]~feeder_combout ;
wire \my_reg[23][13]~q ;
wire \Mux50~17_combout ;
wire \Mux50~18_combout ;
wire \my_reg[28][13]~feeder_combout ;
wire \my_reg[28][13]~q ;
wire \my_reg[24][13]~q ;
wire \Mux50~14_combout ;
wire \Mux50~15_combout ;
wire \my_reg[22][13]~q ;
wire \Mux50~12_combout ;
wire \my_reg[26][13]~q ;
wire \Mux50~13_combout ;
wire \Mux50~16_combout ;
wire \my_reg[24][12]~q ;
wire \my_reg[28][12]~q ;
wire \my_reg[20][12]~q ;
wire \my_reg[16][12]~q ;
wire \Mux19~4_combout ;
wire \Mux19~5_combout ;
wire \my_reg[30][12]~feeder_combout ;
wire \my_reg[30][12]~q ;
wire \my_reg[18][12]~feeder_combout ;
wire \my_reg[18][12]~q ;
wire \Mux19~2_combout ;
wire \Mux19~3_combout ;
wire \Mux19~6_combout ;
wire \my_reg[21][12]~q ;
wire \my_reg[25][12]~feeder_combout ;
wire \my_reg[25][12]~q ;
wire \Mux19~0_combout ;
wire \Mux19~1_combout ;
wire \my_reg[31][12]~feeder_combout ;
wire \my_reg[31][12]~q ;
wire \my_reg[27][12]~q ;
wire \Mux19~7_combout ;
wire \Mux19~8_combout ;
wire \Mux19~9_combout ;
wire \my_reg[1][12]~q ;
wire \Mux19~14_combout ;
wire \Mux19~15_combout ;
wire \my_reg[9][12]~q ;
wire \my_reg[11][12]~q ;
wire \my_reg[8][12]~feeder_combout ;
wire \my_reg[8][12]~q ;
wire \Mux19~12_combout ;
wire \Mux19~13_combout ;
wire \Mux19~16_combout ;
wire \my_reg[12][12]~feeder_combout ;
wire \my_reg[12][12]~q ;
wire \my_reg[13][12]~q ;
wire \Mux19~17_combout ;
wire \my_reg[14][12]~q ;
wire \Mux19~18_combout ;
wire \my_reg[6][12]~feeder_combout ;
wire \my_reg[6][12]~q ;
wire \my_reg[4][12]~q ;
wire \Mux19~10_combout ;
wire \my_reg[7][12]~q ;
wire \Mux19~11_combout ;
wire \Mux19~19_combout ;
wire \my_reg[10][12]~q ;
wire \Mux51~0_combout ;
wire \Mux51~1_combout ;
wire \my_reg[15][12]~q ;
wire \Mux51~7_combout ;
wire \Mux51~8_combout ;
wire \Mux51~2_combout ;
wire \Mux51~3_combout ;
wire \my_reg[2][12]~q ;
wire \my_reg[3][12]~feeder_combout ;
wire \my_reg[3][12]~q ;
wire \Mux51~4_combout ;
wire \Mux51~5_combout ;
wire \Mux51~6_combout ;
wire \Mux51~10_combout ;
wire \my_reg[29][12]~feeder_combout ;
wire \my_reg[29][12]~q ;
wire \Mux51~11_combout ;
wire \my_reg[19][12]~feeder_combout ;
wire \my_reg[19][12]~q ;
wire \Mux51~17_combout ;
wire \Mux51~18_combout ;
wire \Mux51~14_combout ;
wire \Mux51~15_combout ;
wire \my_reg[26][12]~feeder_combout ;
wire \my_reg[26][12]~q ;
wire \Mux51~12_combout ;
wire \Mux51~13_combout ;
wire \Mux51~16_combout ;
wire \my_reg[7][11]~q ;
wire \my_reg[4][11]~q ;
wire \Mux20~12_combout ;
wire \Mux20~13_combout ;
wire \my_reg[1][11]~q ;
wire \my_reg[3][11]~q ;
wire \Mux20~14_combout ;
wire \Mux20~15_combout ;
wire \Mux20~16_combout ;
wire \my_reg[14][11]~q ;
wire \my_reg[13][11]~q ;
wire \Mux20~17_combout ;
wire \Mux20~18_combout ;
wire \my_reg[11][11]~q ;
wire \my_reg[10][11]~q ;
wire \Mux20~10_combout ;
wire \Mux20~11_combout ;
wire \Mux20~19_combout ;
wire \my_reg[31][11]~q ;
wire \my_reg[19][11]~q ;
wire \Mux20~7_combout ;
wire \Mux20~8_combout ;
wire \my_reg[20][11]~q ;
wire \my_reg[28][11]~q ;
wire \my_reg[24][11]~q ;
wire \my_reg[16][11]~q ;
wire \Mux20~4_combout ;
wire \Mux20~5_combout ;
wire \my_reg[30][11]~q ;
wire \my_reg[18][11]~feeder_combout ;
wire \my_reg[18][11]~q ;
wire \Mux20~2_combout ;
wire \Mux20~3_combout ;
wire \Mux20~6_combout ;
wire \my_reg[29][11]~q ;
wire \my_reg[17][11]~q ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \Mux20~9_combout ;
wire \my_reg[12][11]~q ;
wire \Mux52~7_combout ;
wire \my_reg[15][11]~q ;
wire \Mux52~8_combout ;
wire \my_reg[9][11]~feeder_combout ;
wire \my_reg[9][11]~q ;
wire \my_reg[8][11]~q ;
wire \Mux52~2_combout ;
wire \Mux52~3_combout ;
wire \my_reg[2][11]~q ;
wire \Mux52~5_combout ;
wire \Mux52~6_combout ;
wire \my_reg[6][11]~q ;
wire \my_reg[5][11]~q ;
wire \Mux52~0_combout ;
wire \Mux52~1_combout ;
wire \my_reg[27][11]~feeder_combout ;
wire \my_reg[27][11]~q ;
wire \Mux52~17_combout ;
wire \my_reg[23][11]~q ;
wire \Mux52~18_combout ;
wire \my_reg[21][11]~feeder_combout ;
wire \my_reg[21][11]~q ;
wire \my_reg[25][11]~q ;
wire \Mux52~10_combout ;
wire \Mux52~11_combout ;
wire \Mux52~14_combout ;
wire \Mux52~15_combout ;
wire \my_reg[26][11]~q ;
wire \my_reg[22][11]~q ;
wire \Mux52~12_combout ;
wire \Mux52~13_combout ;
wire \Mux52~16_combout ;
wire \my_reg[23][10]~q ;
wire \my_reg[19][10]~feeder_combout ;
wire \my_reg[19][10]~q ;
wire \Mux21~7_combout ;
wire \Mux21~8_combout ;
wire \my_reg[29][10]~q ;
wire \my_reg[21][10]~q ;
wire \Mux21~1_combout ;
wire \my_reg[24][10]~q ;
wire \my_reg[28][10]~q ;
wire \my_reg[20][10]~q ;
wire \my_reg[16][10]~q ;
wire \Mux21~4_combout ;
wire \Mux21~5_combout ;
wire \my_reg[30][10]~q ;
wire \my_reg[18][10]~q ;
wire \Mux21~2_combout ;
wire \Mux21~3_combout ;
wire \Mux21~6_combout ;
wire \Mux21~9_combout ;
wire \my_reg[7][10]~q ;
wire \my_reg[6][10]~q ;
wire \my_reg[4][10]~q ;
wire \my_reg[5][10]~q ;
wire \Mux21~10_combout ;
wire \Mux21~11_combout ;
wire \my_reg[2][10]~q ;
wire \my_reg[1][10]~q ;
wire \my_reg[3][10]~q ;
wire \Mux21~14_combout ;
wire \Mux21~15_combout ;
wire \my_reg[9][10]~feeder_combout ;
wire \my_reg[9][10]~q ;
wire \my_reg[11][10]~q ;
wire \my_reg[8][10]~q ;
wire \Mux21~12_combout ;
wire \Mux21~13_combout ;
wire \Mux21~16_combout ;
wire \my_reg[15][10]~feeder_combout ;
wire \my_reg[15][10]~q ;
wire \my_reg[12][10]~q ;
wire \Mux21~17_combout ;
wire \Mux21~18_combout ;
wire \Mux21~19_combout ;
wire \my_reg[10][10]~feeder_combout ;
wire \my_reg[10][10]~q ;
wire \Mux53~0_combout ;
wire \Mux53~1_combout ;
wire \Mux53~4_combout ;
wire \Mux53~5_combout ;
wire \Mux53~2_combout ;
wire \Mux53~3_combout ;
wire \Mux53~6_combout ;
wire \my_reg[14][10]~feeder_combout ;
wire \my_reg[14][10]~q ;
wire \my_reg[13][10]~feeder_combout ;
wire \my_reg[13][10]~q ;
wire \Mux53~7_combout ;
wire \Mux53~8_combout ;
wire \my_reg[25][10]~q ;
wire \Mux53~10_combout ;
wire \Mux53~11_combout ;
wire \my_reg[31][10]~feeder_combout ;
wire \my_reg[31][10]~q ;
wire \my_reg[27][10]~q ;
wire \Mux53~17_combout ;
wire \Mux53~18_combout ;
wire \Mux53~14_combout ;
wire \Mux53~15_combout ;
wire \my_reg[22][10]~q ;
wire \my_reg[26][10]~q ;
wire \Mux53~12_combout ;
wire \Mux53~13_combout ;
wire \Mux53~16_combout ;
wire \my_reg[25][9]~q ;
wire \my_reg[29][9]~q ;
wire \Mux22~1_combout ;
wire \my_reg[27][9]~feeder_combout ;
wire \my_reg[27][9]~q ;
wire \my_reg[31][9]~q ;
wire \my_reg[19][9]~feeder_combout ;
wire \my_reg[19][9]~q ;
wire \my_reg[23][9]~q ;
wire \Mux22~7_combout ;
wire \Mux22~8_combout ;
wire \my_reg[28][9]~feeder_combout ;
wire \my_reg[28][9]~q ;
wire \my_reg[16][9]~feeder_combout ;
wire \my_reg[16][9]~q ;
wire \Mux22~4_combout ;
wire \Mux22~5_combout ;
wire \my_reg[22][9]~q ;
wire \my_reg[18][9]~feeder_combout ;
wire \my_reg[18][9]~q ;
wire \Mux22~2_combout ;
wire \Mux22~3_combout ;
wire \Mux22~6_combout ;
wire \Mux22~9_combout ;
wire \my_reg[14][9]~q ;
wire \my_reg[13][9]~q ;
wire \Mux22~17_combout ;
wire \Mux22~18_combout ;
wire \my_reg[11][9]~q ;
wire \my_reg[8][9]~q ;
wire \my_reg[10][9]~q ;
wire \Mux22~10_combout ;
wire \Mux22~11_combout ;
wire \my_reg[6][9]~q ;
wire \my_reg[7][9]~q ;
wire \my_reg[4][9]~q ;
wire \Mux22~12_combout ;
wire \Mux22~13_combout ;
wire \my_reg[1][9]~q ;
wire \my_reg[3][9]~q ;
wire \Mux22~14_combout ;
wire \Mux22~15_combout ;
wire \Mux22~16_combout ;
wire \Mux22~19_combout ;
wire \Mux54~2_combout ;
wire \Mux54~3_combout ;
wire \my_reg[2][9]~q ;
wire \Mux54~4_combout ;
wire \Mux54~5_combout ;
wire \Mux54~6_combout ;
wire \my_reg[15][9]~feeder_combout ;
wire \my_reg[15][9]~q ;
wire \my_reg[12][9]~feeder_combout ;
wire \my_reg[12][9]~q ;
wire \Mux54~7_combout ;
wire \Mux54~8_combout ;
wire \my_reg[5][9]~q ;
wire \Mux54~0_combout ;
wire \Mux54~1_combout ;
wire \my_reg[21][9]~feeder_combout ;
wire \my_reg[21][9]~q ;
wire \Mux54~10_combout ;
wire \Mux54~11_combout ;
wire \Mux54~17_combout ;
wire \Mux54~18_combout ;
wire \my_reg[26][9]~q ;
wire \Mux54~12_combout ;
wire \Mux54~13_combout ;
wire \my_reg[24][9]~feeder_combout ;
wire \my_reg[24][9]~q ;
wire \my_reg[20][9]~q ;
wire \Mux54~14_combout ;
wire \Mux54~15_combout ;
wire \Mux54~16_combout ;
wire \my_reg[31][8]~q ;
wire \my_reg[19][8]~feeder_combout ;
wire \my_reg[19][8]~q ;
wire \Mux23~7_combout ;
wire \Mux23~8_combout ;
wire \my_reg[29][8]~q ;
wire \my_reg[25][8]~q ;
wire \Mux23~0_combout ;
wire \Mux23~1_combout ;
wire \my_reg[30][8]~feeder_combout ;
wire \my_reg[30][8]~q ;
wire \my_reg[18][8]~feeder_combout ;
wire \my_reg[18][8]~q ;
wire \Mux23~2_combout ;
wire \Mux23~3_combout ;
wire \my_reg[24][8]~q ;
wire \my_reg[28][8]~q ;
wire \my_reg[20][8]~q ;
wire \my_reg[16][8]~q ;
wire \Mux23~4_combout ;
wire \Mux23~5_combout ;
wire \Mux23~6_combout ;
wire \Mux23~9_combout ;
wire \my_reg[7][8]~q ;
wire \my_reg[6][8]~q ;
wire \my_reg[5][8]~feeder_combout ;
wire \my_reg[5][8]~q ;
wire \Mux23~10_combout ;
wire \Mux23~11_combout ;
wire \my_reg[14][8]~feeder_combout ;
wire \my_reg[14][8]~q ;
wire \my_reg[13][8]~q ;
wire \Mux23~17_combout ;
wire \Mux23~18_combout ;
wire \my_reg[1][8]~q ;
wire \my_reg[3][8]~q ;
wire \Mux23~14_combout ;
wire \Mux23~15_combout ;
wire \my_reg[11][8]~q ;
wire \my_reg[8][8]~q ;
wire \Mux23~12_combout ;
wire \Mux23~13_combout ;
wire \Mux23~16_combout ;
wire \Mux23~19_combout ;
wire \my_reg[12][8]~q ;
wire \Mux55~7_combout ;
wire \my_reg[15][8]~q ;
wire \Mux55~8_combout ;
wire \Mux55~4_combout ;
wire \my_reg[2][8]~q ;
wire \Mux55~5_combout ;
wire \my_reg[4][8]~q ;
wire \Mux55~2_combout ;
wire \Mux55~3_combout ;
wire \Mux55~6_combout ;
wire \my_reg[9][8]~feeder_combout ;
wire \my_reg[9][8]~q ;
wire \my_reg[10][8]~q ;
wire \Mux55~0_combout ;
wire \Mux55~1_combout ;
wire \my_reg[27][8]~feeder_combout ;
wire \my_reg[27][8]~q ;
wire \my_reg[23][8]~q ;
wire \Mux55~17_combout ;
wire \Mux55~18_combout ;
wire \Mux55~14_combout ;
wire \Mux55~15_combout ;
wire \my_reg[26][8]~feeder_combout ;
wire \my_reg[26][8]~q ;
wire \Mux55~12_combout ;
wire \Mux55~13_combout ;
wire \Mux55~16_combout ;
wire \my_reg[17][8]~feeder_combout ;
wire \my_reg[17][8]~q ;
wire \Mux55~10_combout ;
wire \Mux55~11_combout ;
wire \my_reg[27][7]~q ;
wire \my_reg[31][7]~q ;
wire \my_reg[23][7]~q ;
wire \Mux24~7_combout ;
wire \Mux24~8_combout ;
wire \my_reg[25][7]~feeder_combout ;
wire \my_reg[25][7]~q ;
wire \my_reg[29][7]~q ;
wire \my_reg[17][7]~feeder_combout ;
wire \my_reg[17][7]~q ;
wire \my_reg[21][7]~q ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \my_reg[20][7]~feeder_combout ;
wire \my_reg[20][7]~q ;
wire \my_reg[16][7]~q ;
wire \Mux24~4_combout ;
wire \Mux24~5_combout ;
wire \my_reg[22][7]~feeder_combout ;
wire \my_reg[22][7]~q ;
wire \my_reg[26][7]~feeder_combout ;
wire \my_reg[26][7]~q ;
wire \Mux24~2_combout ;
wire \Mux24~3_combout ;
wire \Mux24~6_combout ;
wire \my_reg[9][7]~feeder_combout ;
wire \my_reg[9][7]~q ;
wire \my_reg[11][7]~q ;
wire \my_reg[8][7]~q ;
wire \my_reg[10][7]~q ;
wire \Mux24~10_combout ;
wire \Mux24~11_combout ;
wire \my_reg[4][7]~q ;
wire \Mux24~12_combout ;
wire \my_reg[7][7]~q ;
wire \Mux24~13_combout ;
wire \my_reg[2][7]~q ;
wire \my_reg[3][7]~q ;
wire \Mux24~14_combout ;
wire \Mux24~15_combout ;
wire \Mux24~16_combout ;
wire \my_reg[13][7]~q ;
wire \Mux24~17_combout ;
wire \my_reg[15][7]~feeder_combout ;
wire \my_reg[15][7]~q ;
wire \my_reg[14][7]~q ;
wire \Mux24~18_combout ;
wire \my_reg[12][7]~q ;
wire \Mux56~7_combout ;
wire \Mux56~8_combout ;
wire \Mux56~2_combout ;
wire \Mux56~3_combout ;
wire \my_reg[1][7]~q ;
wire \Mux56~4_combout ;
wire \Mux56~5_combout ;
wire \Mux56~6_combout ;
wire \my_reg[6][7]~q ;
wire \my_reg[5][7]~feeder_combout ;
wire \my_reg[5][7]~q ;
wire \Mux56~0_combout ;
wire \Mux56~1_combout ;
wire \Mux56~17_combout ;
wire \Mux56~18_combout ;
wire \Mux56~10_combout ;
wire \Mux56~11_combout ;
wire \my_reg[18][7]~q ;
wire \Mux56~12_combout ;
wire \my_reg[30][7]~q ;
wire \Mux56~13_combout ;
wire \my_reg[28][7]~q ;
wire \Mux56~14_combout ;
wire \Mux56~15_combout ;
wire \Mux56~16_combout ;
wire \my_reg[21][6]~feeder_combout ;
wire \my_reg[21][6]~q ;
wire \my_reg[25][6]~q ;
wire \Mux25~0_combout ;
wire \my_reg[29][6]~q ;
wire \Mux25~1_combout ;
wire \my_reg[26][6]~feeder_combout ;
wire \my_reg[26][6]~q ;
wire \my_reg[22][6]~feeder_combout ;
wire \my_reg[22][6]~q ;
wire \Mux25~2_combout ;
wire \Mux25~3_combout ;
wire \my_reg[24][6]~feeder_combout ;
wire \my_reg[24][6]~q ;
wire \my_reg[20][6]~q ;
wire \Mux25~4_combout ;
wire \Mux25~5_combout ;
wire \Mux25~6_combout ;
wire \my_reg[31][6]~feeder_combout ;
wire \my_reg[31][6]~q ;
wire \my_reg[23][6]~feeder_combout ;
wire \my_reg[23][6]~q ;
wire \my_reg[27][6]~feeder_combout ;
wire \my_reg[27][6]~q ;
wire \Mux25~7_combout ;
wire \Mux25~8_combout ;
wire \my_reg[14][6]~feeder_combout ;
wire \my_reg[14][6]~q ;
wire \my_reg[15][6]~q ;
wire \my_reg[13][6]~feeder_combout ;
wire \my_reg[13][6]~q ;
wire \Mux25~17_combout ;
wire \Mux25~18_combout ;
wire \my_reg[7][6]~feeder_combout ;
wire \my_reg[7][6]~q ;
wire \my_reg[6][6]~q ;
wire \my_reg[4][6]~feeder_combout ;
wire \my_reg[4][6]~q ;
wire \my_reg[5][6]~q ;
wire \Mux25~10_combout ;
wire \Mux25~11_combout ;
wire \my_reg[10][6]~q ;
wire \my_reg[8][6]~q ;
wire \Mux25~12_combout ;
wire \my_reg[11][6]~q ;
wire \Mux25~13_combout ;
wire \my_reg[3][6]~q ;
wire \Mux25~14_combout ;
wire \Mux25~15_combout ;
wire \Mux25~16_combout ;
wire \my_reg[9][6]~q ;
wire \Mux57~0_combout ;
wire \Mux57~1_combout ;
wire \Mux57~2_combout ;
wire \Mux57~3_combout ;
wire \my_reg[2][6]~q ;
wire \Mux57~4_combout ;
wire \Mux57~5_combout ;
wire \Mux57~6_combout ;
wire \my_reg[12][6]~q ;
wire \Mux57~7_combout ;
wire \Mux57~8_combout ;
wire \Mux57~10_combout ;
wire \Mux57~11_combout ;
wire \my_reg[18][6]~q ;
wire \Mux57~12_combout ;
wire \my_reg[30][6]~q ;
wire \Mux57~13_combout ;
wire \my_reg[16][6]~q ;
wire \Mux57~14_combout ;
wire \my_reg[28][6]~q ;
wire \Mux57~15_combout ;
wire \Mux57~16_combout ;
wire \my_reg[19][6]~q ;
wire \Mux57~17_combout ;
wire \Mux57~18_combout ;
wire \my_reg[11][5]~q ;
wire \my_reg[9][5]~q ;
wire \my_reg[8][5]~q ;
wire \my_reg[10][5]~feeder_combout ;
wire \my_reg[10][5]~q ;
wire \Mux26~10_combout ;
wire \Mux26~11_combout ;
wire \my_reg[2][5]~q ;
wire \my_reg[1][5]~q ;
wire \my_reg[3][5]~q ;
wire \Mux26~14_combout ;
wire \Mux26~15_combout ;
wire \my_reg[7][5]~q ;
wire \my_reg[4][5]~q ;
wire \Mux26~12_combout ;
wire \Mux26~13_combout ;
wire \Mux26~16_combout ;
wire \my_reg[14][5]~feeder_combout ;
wire \my_reg[14][5]~q ;
wire \my_reg[13][5]~q ;
wire \Mux26~17_combout ;
wire \Mux26~18_combout ;
wire \Mux26~19_combout ;
wire \my_reg[27][5]~q ;
wire \my_reg[19][5]~q ;
wire \Mux26~7_combout ;
wire \Mux26~8_combout ;
wire \my_reg[29][5]~q ;
wire \my_reg[21][5]~feeder_combout ;
wire \my_reg[21][5]~q ;
wire \Mux26~0_combout ;
wire \Mux26~1_combout ;
wire \my_reg[28][5]~feeder_combout ;
wire \my_reg[28][5]~q ;
wire \my_reg[20][5]~q ;
wire \my_reg[16][5]~feeder_combout ;
wire \my_reg[16][5]~q ;
wire \Mux26~4_combout ;
wire \Mux26~5_combout ;
wire \my_reg[30][5]~q ;
wire \my_reg[18][5]~q ;
wire \Mux26~2_combout ;
wire \Mux26~3_combout ;
wire \Mux26~6_combout ;
wire \Mux26~9_combout ;
wire \my_reg[6][5]~q ;
wire \my_reg[5][5]~q ;
wire \Mux58~0_combout ;
wire \Mux58~1_combout ;
wire \my_reg[15][5]~q ;
wire \my_reg[12][5]~q ;
wire \Mux58~7_combout ;
wire \Mux58~8_combout ;
wire \Mux58~4_combout ;
wire \Mux58~5_combout ;
wire \Mux58~2_combout ;
wire \Mux58~3_combout ;
wire \Mux58~6_combout ;
wire \Mux58~17_combout ;
wire \my_reg[23][5]~feeder_combout ;
wire \my_reg[23][5]~q ;
wire \my_reg[31][5]~q ;
wire \Mux58~18_combout ;
wire \my_reg[24][5]~feeder_combout ;
wire \my_reg[24][5]~q ;
wire \Mux58~14_combout ;
wire \Mux58~15_combout ;
wire \my_reg[22][5]~feeder_combout ;
wire \my_reg[22][5]~q ;
wire \Mux58~12_combout ;
wire \Mux58~13_combout ;
wire \Mux58~16_combout ;
wire \my_reg[17][5]~q ;
wire \Mux58~10_combout ;
wire \Mux58~11_combout ;
wire \my_reg[29][4]~feeder_combout ;
wire \my_reg[29][4]~q ;
wire \my_reg[21][4]~feeder_combout ;
wire \my_reg[21][4]~q ;
wire \my_reg[25][4]~feeder_combout ;
wire \my_reg[25][4]~q ;
wire \Mux27~0_combout ;
wire \Mux27~1_combout ;
wire \my_reg[31][4]~feeder_combout ;
wire \my_reg[31][4]~q ;
wire \my_reg[23][4]~feeder_combout ;
wire \my_reg[23][4]~q ;
wire \my_reg[19][4]~feeder_combout ;
wire \my_reg[19][4]~q ;
wire \my_reg[27][4]~q ;
wire \Mux27~7_combout ;
wire \Mux27~8_combout ;
wire \my_reg[24][4]~q ;
wire \my_reg[20][4]~q ;
wire \Mux27~4_combout ;
wire \Mux27~5_combout ;
wire \my_reg[26][4]~feeder_combout ;
wire \my_reg[26][4]~q ;
wire \my_reg[18][4]~q ;
wire \Mux27~2_combout ;
wire \Mux27~3_combout ;
wire \Mux27~6_combout ;
wire \my_reg[1][4]~q ;
wire \my_reg[3][4]~q ;
wire \Mux27~14_combout ;
wire \Mux27~15_combout ;
wire \my_reg[9][4]~feeder_combout ;
wire \my_reg[9][4]~q ;
wire \my_reg[8][4]~q ;
wire \my_reg[10][4]~q ;
wire \Mux27~12_combout ;
wire \Mux27~13_combout ;
wire \Mux27~16_combout ;
wire \my_reg[15][4]~q ;
wire \my_reg[14][4]~feeder_combout ;
wire \my_reg[14][4]~q ;
wire \my_reg[13][4]~q ;
wire \Mux27~17_combout ;
wire \Mux27~18_combout ;
wire \my_reg[7][4]~feeder_combout ;
wire \my_reg[7][4]~q ;
wire \my_reg[6][4]~q ;
wire \my_reg[4][4]~feeder_combout ;
wire \my_reg[4][4]~q ;
wire \my_reg[5][4]~q ;
wire \Mux27~10_combout ;
wire \Mux27~11_combout ;
wire \my_reg[11][4]~q ;
wire \Mux59~0_combout ;
wire \Mux59~1_combout ;
wire \my_reg[12][4]~q ;
wire \Mux59~7_combout ;
wire \Mux59~8_combout ;
wire \my_reg[2][4]~q ;
wire \Mux59~4_combout ;
wire \Mux59~5_combout ;
wire \Mux59~2_combout ;
wire \Mux59~3_combout ;
wire \Mux59~6_combout ;
wire \Mux59~17_combout ;
wire \Mux59~18_combout ;
wire \my_reg[28][4]~q ;
wire \my_reg[16][4]~q ;
wire \Mux59~14_combout ;
wire \Mux59~15_combout ;
wire \my_reg[22][4]~feeder_combout ;
wire \my_reg[22][4]~q ;
wire \my_reg[30][4]~q ;
wire \Mux59~12_combout ;
wire \Mux59~13_combout ;
wire \Mux59~16_combout ;
wire \my_reg[17][4]~feeder_combout ;
wire \my_reg[17][4]~q ;
wire \Mux59~10_combout ;
wire \Mux59~11_combout ;
wire \my_reg[14][3]~feeder_combout ;
wire \my_reg[14][3]~q ;
wire \my_reg[12][3]~feeder_combout ;
wire \my_reg[12][3]~q ;
wire \my_reg[13][3]~q ;
wire \Mux28~17_combout ;
wire \my_reg[15][3]~q ;
wire \Mux28~18_combout ;
wire \my_reg[7][3]~q ;
wire \my_reg[4][3]~q ;
wire \Mux28~12_combout ;
wire \Mux28~13_combout ;
wire \my_reg[2][3]~q ;
wire \my_reg[3][3]~feeder_combout ;
wire \my_reg[3][3]~q ;
wire \Mux28~14_combout ;
wire \Mux28~15_combout ;
wire \Mux28~16_combout ;
wire \my_reg[11][3]~q ;
wire \my_reg[9][3]~q ;
wire \my_reg[8][3]~q ;
wire \my_reg[10][3]~q ;
wire \Mux28~10_combout ;
wire \Mux28~11_combout ;
wire \Mux28~19_combout ;
wire \my_reg[29][3]~q ;
wire \my_reg[17][3]~q ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \my_reg[31][3]~feeder_combout ;
wire \my_reg[31][3]~q ;
wire \my_reg[27][3]~q ;
wire \my_reg[23][3]~q ;
wire \Mux28~7_combout ;
wire \Mux28~8_combout ;
wire \my_reg[30][3]~q ;
wire \my_reg[18][3]~feeder_combout ;
wire \my_reg[18][3]~q ;
wire \Mux28~2_combout ;
wire \Mux28~3_combout ;
wire \Mux28~6_combout ;
wire \Mux28~9_combout ;
wire \my_reg[19][3]~feeder_combout ;
wire \my_reg[19][3]~q ;
wire \Mux60~7_combout ;
wire \Mux60~8_combout ;
wire \my_reg[21][3]~feeder_combout ;
wire \my_reg[21][3]~q ;
wire \my_reg[25][3]~feeder_combout ;
wire \my_reg[25][3]~q ;
wire \Mux60~0_combout ;
wire \Mux60~1_combout ;
wire \my_reg[26][3]~feeder_combout ;
wire \my_reg[26][3]~q ;
wire \my_reg[22][3]~q ;
wire \Mux60~2_combout ;
wire \Mux60~3_combout ;
wire \my_reg[28][3]~feeder_combout ;
wire \my_reg[28][3]~q ;
wire \my_reg[20][3]~feeder_combout ;
wire \my_reg[20][3]~q ;
wire \Mux60~4_combout ;
wire \Mux60~5_combout ;
wire \Mux60~6_combout ;
wire \my_reg[6][3]~q ;
wire \my_reg[5][3]~q ;
wire \Mux60~10_combout ;
wire \Mux60~11_combout ;
wire \Mux60~17_combout ;
wire \Mux60~18_combout ;
wire \my_reg[1][3]~q ;
wire \Mux60~14_combout ;
wire \Mux60~15_combout ;
wire \Mux60~12_combout ;
wire \Mux60~13_combout ;
wire \Mux60~16_combout ;
wire \my_reg[31][2]~feeder_combout ;
wire \my_reg[31][2]~q ;
wire \my_reg[23][2]~feeder_combout ;
wire \my_reg[23][2]~q ;
wire \my_reg[19][2]~feeder_combout ;
wire \my_reg[19][2]~q ;
wire \Mux29~7_combout ;
wire \Mux29~8_combout ;
wire \my_reg[21][2]~q ;
wire \my_reg[25][2]~q ;
wire \Mux29~0_combout ;
wire \my_reg[29][2]~feeder_combout ;
wire \my_reg[29][2]~q ;
wire \Mux29~1_combout ;
wire \my_reg[24][2]~feeder_combout ;
wire \my_reg[24][2]~q ;
wire \my_reg[16][2]~q ;
wire \Mux29~4_combout ;
wire \Mux29~5_combout ;
wire \my_reg[30][2]~q ;
wire \my_reg[18][2]~q ;
wire \Mux29~2_combout ;
wire \Mux29~3_combout ;
wire \Mux29~6_combout ;
wire \my_reg[14][2]~feeder_combout ;
wire \my_reg[14][2]~q ;
wire \my_reg[15][2]~q ;
wire \my_reg[13][2]~feeder_combout ;
wire \my_reg[13][2]~q ;
wire \Mux29~17_combout ;
wire \Mux29~18_combout ;
wire \my_reg[6][2]~feeder_combout ;
wire \my_reg[6][2]~q ;
wire \my_reg[7][2]~feeder_combout ;
wire \my_reg[7][2]~q ;
wire \my_reg[4][2]~feeder_combout ;
wire \my_reg[4][2]~q ;
wire \my_reg[5][2]~q ;
wire \Mux29~10_combout ;
wire \Mux29~11_combout ;
wire \my_reg[9][2]~feeder_combout ;
wire \my_reg[9][2]~q ;
wire \my_reg[8][2]~feeder_combout ;
wire \my_reg[8][2]~q ;
wire \Mux29~12_combout ;
wire \Mux29~13_combout ;
wire \my_reg[3][2]~feeder_combout ;
wire \my_reg[3][2]~q ;
wire \Mux29~14_combout ;
wire \my_reg[2][2]~feeder_combout ;
wire \my_reg[2][2]~q ;
wire \Mux29~15_combout ;
wire \Mux29~16_combout ;
wire \my_reg[11][2]~feeder_combout ;
wire \my_reg[11][2]~q ;
wire \Mux61~0_combout ;
wire \Mux61~1_combout ;
wire \my_reg[12][2]~feeder_combout ;
wire \my_reg[12][2]~q ;
wire \Mux61~7_combout ;
wire \Mux61~8_combout ;
wire \my_reg[1][2]~q ;
wire \Mux61~4_combout ;
wire \Mux61~5_combout ;
wire \Mux61~2_combout ;
wire \Mux61~3_combout ;
wire \Mux61~6_combout ;
wire \my_reg[17][2]~feeder_combout ;
wire \my_reg[17][2]~q ;
wire \Mux61~10_combout ;
wire \Mux61~11_combout ;
wire \my_reg[27][2]~feeder_combout ;
wire \my_reg[27][2]~q ;
wire \Mux61~17_combout ;
wire \Mux61~18_combout ;
wire \my_reg[28][2]~q ;
wire \Mux61~14_combout ;
wire \Mux61~15_combout ;
wire \my_reg[22][2]~feeder_combout ;
wire \my_reg[22][2]~q ;
wire \my_reg[26][2]~feeder_combout ;
wire \my_reg[26][2]~q ;
wire \Mux61~12_combout ;
wire \Mux61~13_combout ;
wire \Mux61~16_combout ;
wire \my_reg[17][1]~feeder_combout ;
wire \my_reg[17][1]~q ;
wire \Mux62~0_combout ;
wire \Mux62~1_combout ;
wire \my_reg[19][1]~feeder_combout ;
wire \my_reg[19][1]~q ;
wire \Mux62~7_combout ;
wire \Mux62~8_combout ;
wire \my_reg[28][1]~feeder_combout ;
wire \my_reg[28][1]~q ;
wire \Mux62~4_combout ;
wire \Mux62~5_combout ;
wire \my_reg[26][1]~q ;
wire \Mux62~2_combout ;
wire \Mux62~3_combout ;
wire \Mux62~6_combout ;
wire \Mux62~10_combout ;
wire \Mux62~11_combout ;
wire \my_reg[12][1]~feeder_combout ;
wire \my_reg[12][1]~q ;
wire \Mux62~19_combout ;
wire \Mux62~20_combout ;
wire \Mux62~15_combout ;
wire \Mux62~16_combout ;
wire \Mux62~17_combout ;
wire \Mux62~12_combout ;
wire \Mux62~13_combout ;
wire \Mux62~18_combout ;
wire \my_reg[22][0]~feeder_combout ;
wire \my_reg[22][0]~q ;
wire \Mux31~2_combout ;
wire \Mux31~3_combout ;
wire \my_reg[28][0]~feeder_combout ;
wire \my_reg[28][0]~q ;
wire \Mux31~4_combout ;
wire \Mux31~5_combout ;
wire \Mux31~6_combout ;
wire \my_reg[17][0]~q ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \my_reg[19][0]~feeder_combout ;
wire \my_reg[19][0]~q ;
wire \Mux31~7_combout ;
wire \Mux31~8_combout ;
wire \Mux31~17_combout ;
wire \Mux31~18_combout ;
wire \my_reg[8][0]~q ;
wire \Mux31~12_combout ;
wire \Mux31~13_combout ;
wire \Mux31~14_combout ;
wire \Mux31~15_combout ;
wire \Mux31~16_combout ;
wire \Mux31~10_combout ;
wire \Mux31~11_combout ;


// Location: FF_X61_Y35_N29
dffeas \my_reg[4][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][0] .is_wysiwyg = "true";
defparam \my_reg[4][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N14
cycloneive_lcell_comb \Mux63~12 (
// Equation(s):
// \Mux63~12_combout  = (instr_16 & ((instr_17) # ((\my_reg[5][0]~q )))) # (!instr_16 & (!instr_17 & ((\my_reg[4][0]~q ))))

	.dataa(instr_16),
	.datab(instr_17),
	.datac(\my_reg[5][0]~q ),
	.datad(\my_reg[4][0]~q ),
	.cin(gnd),
	.combout(\Mux63~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~12 .lut_mask = 16'hB9A8;
defparam \Mux63~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N0
cycloneive_lcell_comb \Mux63~16 (
// Equation(s):
// \Mux63~16_combout  = (instr_16 & ((instr_17 & ((\my_reg[3][0]~q ))) # (!instr_17 & (\my_reg[1][0]~q ))))

	.dataa(\my_reg[1][0]~q ),
	.datab(instr_17),
	.datac(\my_reg[3][0]~q ),
	.datad(instr_16),
	.cin(gnd),
	.combout(\Mux63~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~16 .lut_mask = 16'hE200;
defparam \Mux63~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N5
dffeas \my_reg[22][1] (
	.clk(CLK),
	.d(\my_reg[22][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][1] .is_wysiwyg = "true";
defparam \my_reg[22][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N23
dffeas \my_reg[24][1] (
	.clk(CLK),
	.d(\my_reg[24][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][1] .is_wysiwyg = "true";
defparam \my_reg[24][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N12
cycloneive_lcell_comb \Mux0~4 (
// Equation(s):
// \Mux0~4_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[24][31]~q )) # (!dcifimemload_24 & ((\my_reg[16][31]~q )))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[24][31]~q ),
	.datac(\my_reg[16][31]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~4 .lut_mask = 16'hEE50;
defparam \Mux0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y42_N13
dffeas \my_reg[10][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][31] .is_wysiwyg = "true";
defparam \my_reg[10][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N21
dffeas \my_reg[5][31] (
	.clk(CLK),
	.d(\my_reg[5][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][31] .is_wysiwyg = "true";
defparam \my_reg[5][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N12
cycloneive_lcell_comb \Mux32~2 (
// Equation(s):
// \Mux32~2_combout  = (dcifimemload_17 & (((\my_reg[10][31]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\my_reg[8][31]~q  & ((!dcifimemload_16))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[8][31]~q ),
	.datac(\my_reg[10][31]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux32~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~2 .lut_mask = 16'hAAE4;
defparam \Mux32~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y38_N13
dffeas \my_reg[10][30] (
	.clk(CLK),
	.d(\my_reg[10][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][30] .is_wysiwyg = "true";
defparam \my_reg[10][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N9
dffeas \my_reg[17][29] (
	.clk(CLK),
	.d(\my_reg[17][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][29] .is_wysiwyg = "true";
defparam \my_reg[17][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N9
dffeas \my_reg[21][28] (
	.clk(CLK),
	.d(\my_reg[21][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][28] .is_wysiwyg = "true";
defparam \my_reg[21][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N3
dffeas \my_reg[12][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][28] .is_wysiwyg = "true";
defparam \my_reg[12][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N2
cycloneive_lcell_comb \Mux3~17 (
// Equation(s):
// \Mux3~17_combout  = (dcifimemload_21 & ((\my_reg[13][28]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][28]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[13][28]~q ),
	.datac(\my_reg[12][28]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux3~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~17 .lut_mask = 16'hAAD8;
defparam \Mux3~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N30
cycloneive_lcell_comb \Mux5~4 (
// Equation(s):
// \Mux5~4_combout  = (dcifimemload_23 & ((\my_reg[20][26]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[16][26]~q  & !dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[20][26]~q ),
	.datac(\my_reg[16][26]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~4 .lut_mask = 16'hAAD8;
defparam \Mux5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N11
dffeas \my_reg[23][26] (
	.clk(CLK),
	.d(\my_reg[23][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][26] .is_wysiwyg = "true";
defparam \my_reg[23][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N27
dffeas \my_reg[2][26] (
	.clk(CLK),
	.d(\my_reg[2][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][26] .is_wysiwyg = "true";
defparam \my_reg[2][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N5
dffeas \my_reg[1][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][25] .is_wysiwyg = "true";
defparam \my_reg[1][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N4
cycloneive_lcell_comb \Mux6~14 (
// Equation(s):
// \Mux6~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\my_reg[3][25]~q )) # (!dcifimemload_22 & ((\my_reg[1][25]~q )))))

	.dataa(\my_reg[3][25]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[1][25]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux6~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~14 .lut_mask = 16'h88C0;
defparam \Mux6~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N22
cycloneive_lcell_comb \Mux8~10 (
// Equation(s):
// \Mux8~10_combout  = (dcifimemload_22 & ((\my_reg[10][23]~q ) # ((dcifimemload_21)))) # (!dcifimemload_22 & (((!dcifimemload_21 & \my_reg[8][23]~q ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[10][23]~q ),
	.datac(dcifimemload_21),
	.datad(\my_reg[8][23]~q ),
	.cin(gnd),
	.combout(\Mux8~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~10 .lut_mask = 16'hADA8;
defparam \Mux8~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N27
dffeas \my_reg[13][23] (
	.clk(CLK),
	.d(\my_reg[13][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][23] .is_wysiwyg = "true";
defparam \my_reg[13][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y42_N27
dffeas \my_reg[5][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][22] .is_wysiwyg = "true";
defparam \my_reg[5][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N3
dffeas \my_reg[3][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][22] .is_wysiwyg = "true";
defparam \my_reg[3][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N26
cycloneive_lcell_comb \Mux41~2 (
// Equation(s):
// \Mux41~2_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][22]~q ))) # (!dcifimemload_16 & (\my_reg[4][22]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[4][22]~q ),
	.datac(\my_reg[5][22]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux41~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~2 .lut_mask = 16'hFA44;
defparam \Mux41~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N12
cycloneive_lcell_comb \Mux41~4 (
// Equation(s):
// \Mux41~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][22]~q ))) # (!dcifimemload_17 & (\my_reg[1][22]~q ))))

	.dataa(\my_reg[1][22]~q ),
	.datab(\my_reg[3][22]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux41~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~4 .lut_mask = 16'hCA00;
defparam \Mux41~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y39_N1
dffeas \my_reg[1][21] (
	.clk(CLK),
	.d(wdat12),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][21] .is_wysiwyg = "true";
defparam \my_reg[1][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N12
cycloneive_lcell_comb \Mux10~14 (
// Equation(s):
// \Mux10~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][21]~q ))) # (!dcifimemload_22 & (\my_reg[1][21]~q ))))

	.dataa(\my_reg[1][21]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[3][21]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux10~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~14 .lut_mask = 16'hC088;
defparam \Mux10~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N7
dffeas \my_reg[12][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][21] .is_wysiwyg = "true";
defparam \my_reg[12][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N6
cycloneive_lcell_comb \Mux10~17 (
// Equation(s):
// \Mux10~17_combout  = (dcifimemload_21 & ((\my_reg[13][21]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][21]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[13][21]~q ),
	.datac(\my_reg[12][21]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux10~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~17 .lut_mask = 16'hAAD8;
defparam \Mux10~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N30
cycloneive_lcell_comb \Mux42~2 (
// Equation(s):
// \Mux42~2_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[10][21]~q ))) # (!dcifimemload_17 & (\my_reg[8][21]~q ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[8][21]~q ),
	.datac(\my_reg[10][21]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux42~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~2 .lut_mask = 16'hFA44;
defparam \Mux42~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N4
cycloneive_lcell_comb \Mux11~12 (
// Equation(s):
// \Mux11~12_combout  = (dcifimemload_22 & ((\my_reg[10][20]~q ) # ((dcifimemload_21)))) # (!dcifimemload_22 & (((\my_reg[8][20]~q  & !dcifimemload_21))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[10][20]~q ),
	.datac(\my_reg[8][20]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux11~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~12 .lut_mask = 16'hAAD8;
defparam \Mux11~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N22
cycloneive_lcell_comb \Mux11~13 (
// Equation(s):
// \Mux11~13_combout  = (\Mux11~12_combout  & (((\my_reg[11][20]~q ) # (!dcifimemload_21)))) # (!\Mux11~12_combout  & (\my_reg[9][20]~q  & ((dcifimemload_21))))

	.dataa(\my_reg[9][20]~q ),
	.datab(\Mux11~12_combout ),
	.datac(\my_reg[11][20]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux11~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~13 .lut_mask = 16'hE2CC;
defparam \Mux11~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N15
dffeas \my_reg[27][19] (
	.clk(CLK),
	.d(\my_reg[27][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][19] .is_wysiwyg = "true";
defparam \my_reg[27][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y32_N27
dffeas \my_reg[5][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][18] .is_wysiwyg = "true";
defparam \my_reg[5][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N26
cycloneive_lcell_comb \Mux45~2 (
// Equation(s):
// \Mux45~2_combout  = (dcifimemload_16 & (((\my_reg[5][18]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[4][18]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[4][18]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[5][18]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux45~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~2 .lut_mask = 16'hCCE2;
defparam \Mux45~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y31_N13
dffeas \my_reg[20][17] (
	.clk(CLK),
	.d(\my_reg[20][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][17] .is_wysiwyg = "true";
defparam \my_reg[20][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N8
cycloneive_lcell_comb \Mux15~2 (
// Equation(s):
// \Mux15~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[22][16]~q )) # (!dcifimemload_23 & ((\my_reg[18][16]~q )))))

	.dataa(\my_reg[22][16]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[18][16]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux15~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~2 .lut_mask = 16'hEE30;
defparam \Mux15~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N13
dffeas \my_reg[30][16] (
	.clk(CLK),
	.d(\my_reg[30][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][16] .is_wysiwyg = "true";
defparam \my_reg[30][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N2
cycloneive_lcell_comb \Mux15~3 (
// Equation(s):
// \Mux15~3_combout  = (\Mux15~2_combout  & ((\my_reg[30][16]~q ) # ((!dcifimemload_24)))) # (!\Mux15~2_combout  & (((\my_reg[26][16]~q  & dcifimemload_24))))

	.dataa(\my_reg[30][16]~q ),
	.datab(\my_reg[26][16]~q ),
	.datac(\Mux15~2_combout ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux15~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~3 .lut_mask = 16'hACF0;
defparam \Mux15~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y30_N23
dffeas \my_reg[20][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][15] .is_wysiwyg = "true";
defparam \my_reg[20][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N31
dffeas \my_reg[27][15] (
	.clk(CLK),
	.d(\my_reg[27][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][15] .is_wysiwyg = "true";
defparam \my_reg[27][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N22
cycloneive_lcell_comb \Mux48~14 (
// Equation(s):
// \Mux48~14_combout  = (dcifimemload_18 & ((dcifimemload_19) # ((\my_reg[20][15]~q )))) # (!dcifimemload_18 & (!dcifimemload_19 & ((\my_reg[16][15]~q ))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\my_reg[20][15]~q ),
	.datad(\my_reg[16][15]~q ),
	.cin(gnd),
	.combout(\Mux48~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~14 .lut_mask = 16'hB9A8;
defparam \Mux48~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N7
dffeas \my_reg[17][14] (
	.clk(CLK),
	.d(\my_reg[17][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][14] .is_wysiwyg = "true";
defparam \my_reg[17][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N26
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (dcifimemload_24 & (((\my_reg[25][14]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\my_reg[17][14]~q  & ((!dcifimemload_23))))

	.dataa(\my_reg[17][14]~q ),
	.datab(\my_reg[25][14]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hF0CA;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y31_N31
dffeas \my_reg[24][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][14] .is_wysiwyg = "true";
defparam \my_reg[24][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N19
dffeas \my_reg[5][14] (
	.clk(CLK),
	.d(\my_reg[5][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][14] .is_wysiwyg = "true";
defparam \my_reg[5][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N30
cycloneive_lcell_comb \Mux49~14 (
// Equation(s):
// \Mux49~14_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[24][14]~q ))) # (!dcifimemload_19 & (\my_reg[16][14]~q ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[16][14]~q ),
	.datac(\my_reg[24][14]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux49~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~14 .lut_mask = 16'hFA44;
defparam \Mux49~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N9
dffeas \my_reg[18][13] (
	.clk(CLK),
	.d(\my_reg[18][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][13] .is_wysiwyg = "true";
defparam \my_reg[18][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N22
cycloneive_lcell_comb \Mux18~2 (
// Equation(s):
// \Mux18~2_combout  = (dcifimemload_24 & ((\my_reg[26][13]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\my_reg[18][13]~q  & !dcifimemload_23))))

	.dataa(\my_reg[26][13]~q ),
	.datab(\my_reg[18][13]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~2 .lut_mask = 16'hF0AC;
defparam \Mux18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y42_N5
dffeas \my_reg[30][13] (
	.clk(CLK),
	.d(\my_reg[30][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][13] .is_wysiwyg = "true";
defparam \my_reg[30][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N26
cycloneive_lcell_comb \Mux18~3 (
// Equation(s):
// \Mux18~3_combout  = (\Mux18~2_combout  & (((\my_reg[30][13]~q ) # (!dcifimemload_23)))) # (!\Mux18~2_combout  & (\my_reg[22][13]~q  & ((dcifimemload_23))))

	.dataa(\my_reg[22][13]~q ),
	.datab(\my_reg[30][13]~q ),
	.datac(\Mux18~2_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~3 .lut_mask = 16'hCAF0;
defparam \Mux18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y39_N15
dffeas \my_reg[1][13] (
	.clk(CLK),
	.d(\my_reg[1][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][13] .is_wysiwyg = "true";
defparam \my_reg[1][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N28
cycloneive_lcell_comb \Mux18~14 (
// Equation(s):
// \Mux18~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][13]~q ))) # (!dcifimemload_22 & (\my_reg[1][13]~q ))))

	.dataa(\my_reg[1][13]~q ),
	.datab(\my_reg[3][13]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux18~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~14 .lut_mask = 16'hC0A0;
defparam \Mux18~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N11
dffeas \my_reg[12][13] (
	.clk(CLK),
	.d(\my_reg[12][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][13] .is_wysiwyg = "true";
defparam \my_reg[12][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N23
dffeas \my_reg[17][12] (
	.clk(CLK),
	.d(\my_reg[17][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][12] .is_wysiwyg = "true";
defparam \my_reg[17][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N31
dffeas \my_reg[22][12] (
	.clk(CLK),
	.d(\my_reg[22][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][12] .is_wysiwyg = "true";
defparam \my_reg[22][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N17
dffeas \my_reg[23][12] (
	.clk(CLK),
	.d(\my_reg[23][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][12] .is_wysiwyg = "true";
defparam \my_reg[23][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N31
dffeas \my_reg[5][12] (
	.clk(CLK),
	.d(\my_reg[5][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][12] .is_wysiwyg = "true";
defparam \my_reg[5][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N6
cycloneive_lcell_comb \Mux52~4 (
// Equation(s):
// \Mux52~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\my_reg[3][11]~q )) # (!dcifimemload_17 & ((\my_reg[1][11]~q )))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[3][11]~q ),
	.datac(\my_reg[1][11]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux52~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~4 .lut_mask = 16'hD800;
defparam \Mux52~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N15
dffeas \my_reg[17][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][10] .is_wysiwyg = "true";
defparam \my_reg[17][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N14
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[25][10]~q )) # (!dcifimemload_24 & ((\my_reg[17][10]~q )))))

	.dataa(\my_reg[25][10]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[17][10]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hEE30;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N29
dffeas \my_reg[17][9] (
	.clk(CLK),
	.d(\my_reg[17][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][9] .is_wysiwyg = "true";
defparam \my_reg[17][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N6
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (dcifimemload_23 & (((\my_reg[21][9]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\my_reg[17][9]~q  & ((!dcifimemload_24))))

	.dataa(\my_reg[17][9]~q ),
	.datab(\my_reg[21][9]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hF0CA;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N13
dffeas \my_reg[30][9] (
	.clk(CLK),
	.d(\my_reg[30][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][9] .is_wysiwyg = "true";
defparam \my_reg[30][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N31
dffeas \my_reg[9][9] (
	.clk(CLK),
	.d(\my_reg[9][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][9] .is_wysiwyg = "true";
defparam \my_reg[9][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N27
dffeas \my_reg[21][8] (
	.clk(CLK),
	.d(\my_reg[21][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][8] .is_wysiwyg = "true";
defparam \my_reg[21][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y43_N11
dffeas \my_reg[22][8] (
	.clk(CLK),
	.d(\my_reg[22][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][8] .is_wysiwyg = "true";
defparam \my_reg[22][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y31_N27
dffeas \my_reg[24][7] (
	.clk(CLK),
	.d(\my_reg[24][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][7] .is_wysiwyg = "true";
defparam \my_reg[24][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y36_N13
dffeas \my_reg[19][7] (
	.clk(CLK),
	.d(\my_reg[19][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][7] .is_wysiwyg = "true";
defparam \my_reg[19][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N27
dffeas \my_reg[17][6] (
	.clk(CLK),
	.d(\my_reg[17][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][6] .is_wysiwyg = "true";
defparam \my_reg[17][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N17
dffeas \my_reg[1][6] (
	.clk(CLK),
	.d(\my_reg[1][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][6] .is_wysiwyg = "true";
defparam \my_reg[1][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N27
dffeas \my_reg[25][5] (
	.clk(CLK),
	.d(\my_reg[25][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][5] .is_wysiwyg = "true";
defparam \my_reg[25][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y43_N3
dffeas \my_reg[26][5] (
	.clk(CLK),
	.d(\my_reg[26][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][5] .is_wysiwyg = "true";
defparam \my_reg[26][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N7
dffeas \my_reg[24][3] (
	.clk(CLK),
	.d(\my_reg[24][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][3] .is_wysiwyg = "true";
defparam \my_reg[24][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N5
dffeas \my_reg[16][3] (
	.clk(CLK),
	.d(\my_reg[16][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][3] .is_wysiwyg = "true";
defparam \my_reg[16][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N2
cycloneive_lcell_comb \Mux28~4 (
// Equation(s):
// \Mux28~4_combout  = (dcifimemload_24 & ((\my_reg[24][3]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\my_reg[16][3]~q  & !dcifimemload_23))))

	.dataa(\my_reg[24][3]~q ),
	.datab(\my_reg[16][3]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~4 .lut_mask = 16'hF0AC;
defparam \Mux28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N6
cycloneive_lcell_comb \Mux28~5 (
// Equation(s):
// \Mux28~5_combout  = (dcifimemload_23 & ((\Mux28~4_combout  & (\my_reg[28][3]~q )) # (!\Mux28~4_combout  & ((\my_reg[20][3]~q ))))) # (!dcifimemload_23 & (((\Mux28~4_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[28][3]~q ),
	.datac(\my_reg[20][3]~q ),
	.datad(\Mux28~4_combout ),
	.cin(gnd),
	.combout(\Mux28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~5 .lut_mask = 16'hDDA0;
defparam \Mux28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y31_N31
dffeas \my_reg[20][2] (
	.clk(CLK),
	.d(\my_reg[20][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][2] .is_wysiwyg = "true";
defparam \my_reg[20][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N21
dffeas \my_reg[10][2] (
	.clk(CLK),
	.d(\my_reg[10][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][2] .is_wysiwyg = "true";
defparam \my_reg[10][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N26
cycloneive_lcell_comb \Mux62~14 (
// Equation(s):
// \Mux62~14_combout  = (instr_16 & ((instr_17 & ((\my_reg[3][1]~q ))) # (!instr_17 & (\my_reg[1][1]~q ))))

	.dataa(\my_reg[1][1]~q ),
	.datab(\my_reg[3][1]~q ),
	.datac(instr_16),
	.datad(instr_17),
	.cin(gnd),
	.combout(\Mux62~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~14 .lut_mask = 16'hC0A0;
defparam \Mux62~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N22
cycloneive_lcell_comb \Decoder0~50 (
// Equation(s):
// \Decoder0~50_combout  = (\wsel~1_combout  & (!\wsel~0_combout  & cuifRegWEN1))

	.dataa(wsel1),
	.datab(gnd),
	.datac(wsel),
	.datad(cuifRegWEN),
	.cin(gnd),
	.combout(\Decoder0~50_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~50 .lut_mask = 16'h0A00;
defparam \Decoder0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N22
cycloneive_lcell_comb \my_reg[24][1]~feeder (
// Equation(s):
// \my_reg[24][1]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\my_reg[24][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[24][1]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[24][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N4
cycloneive_lcell_comb \my_reg[22][1]~feeder (
// Equation(s):
// \my_reg[22][1]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\my_reg[22][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[22][1]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[22][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N20
cycloneive_lcell_comb \my_reg[5][31]~feeder (
// Equation(s):
// \my_reg[5][31]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat2),
	.cin(gnd),
	.combout(\my_reg[5][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[5][31]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[5][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N12
cycloneive_lcell_comb \my_reg[10][30]~feeder (
// Equation(s):
// \my_reg[10][30]~feeder_combout  = \wdat~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat3),
	.cin(gnd),
	.combout(\my_reg[10][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[10][30]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[10][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N8
cycloneive_lcell_comb \my_reg[17][29]~feeder (
// Equation(s):
// \my_reg[17][29]~feeder_combout  = \wdat~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat4),
	.cin(gnd),
	.combout(\my_reg[17][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[17][29]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[17][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N8
cycloneive_lcell_comb \my_reg[21][28]~feeder (
// Equation(s):
// \my_reg[21][28]~feeder_combout  = \wdat~11_combout 

	.dataa(wdat5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[21][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][28]~feeder .lut_mask = 16'hAAAA;
defparam \my_reg[21][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N10
cycloneive_lcell_comb \my_reg[23][26]~feeder (
// Equation(s):
// \my_reg[23][26]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat7),
	.cin(gnd),
	.combout(\my_reg[23][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[23][26]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[23][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N26
cycloneive_lcell_comb \my_reg[2][26]~feeder (
// Equation(s):
// \my_reg[2][26]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat7),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[2][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[2][26]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[2][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N26
cycloneive_lcell_comb \my_reg[13][23]~feeder (
// Equation(s):
// \my_reg[13][23]~feeder_combout  = \wdat~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat10),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[13][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[13][23]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[13][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N14
cycloneive_lcell_comb \my_reg[27][19]~feeder (
// Equation(s):
// \my_reg[27][19]~feeder_combout  = \wdat~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat14),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[27][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[27][19]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[27][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N12
cycloneive_lcell_comb \my_reg[20][17]~feeder (
// Equation(s):
// \my_reg[20][17]~feeder_combout  = \wdat~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat16),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[20][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[20][17]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[20][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N12
cycloneive_lcell_comb \my_reg[30][16]~feeder (
// Equation(s):
// \my_reg[30][16]~feeder_combout  = \wdat~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat17),
	.cin(gnd),
	.combout(\my_reg[30][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[30][16]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[30][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N30
cycloneive_lcell_comb \my_reg[27][15]~feeder (
// Equation(s):
// \my_reg[27][15]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat18),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[27][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[27][15]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[27][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N6
cycloneive_lcell_comb \my_reg[17][14]~feeder (
// Equation(s):
// \my_reg[17][14]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat19),
	.cin(gnd),
	.combout(\my_reg[17][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[17][14]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[17][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N18
cycloneive_lcell_comb \my_reg[5][14]~feeder (
// Equation(s):
// \my_reg[5][14]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat19),
	.cin(gnd),
	.combout(\my_reg[5][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[5][14]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[5][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N14
cycloneive_lcell_comb \my_reg[1][13]~feeder (
// Equation(s):
// \my_reg[1][13]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat20),
	.cin(gnd),
	.combout(\my_reg[1][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[1][13]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[1][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N10
cycloneive_lcell_comb \my_reg[12][13]~feeder (
// Equation(s):
// \my_reg[12][13]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat20),
	.cin(gnd),
	.combout(\my_reg[12][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[12][13]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[12][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N4
cycloneive_lcell_comb \my_reg[30][13]~feeder (
// Equation(s):
// \my_reg[30][13]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat20),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[30][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[30][13]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[30][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N8
cycloneive_lcell_comb \my_reg[18][13]~feeder (
// Equation(s):
// \my_reg[18][13]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat20),
	.cin(gnd),
	.combout(\my_reg[18][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[18][13]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[18][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N30
cycloneive_lcell_comb \my_reg[5][12]~feeder (
// Equation(s):
// \my_reg[5][12]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat21),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[5][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[5][12]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[5][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N30
cycloneive_lcell_comb \my_reg[22][12]~feeder (
// Equation(s):
// \my_reg[22][12]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat21),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[22][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[22][12]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[22][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N22
cycloneive_lcell_comb \my_reg[17][12]~feeder (
// Equation(s):
// \my_reg[17][12]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat21),
	.cin(gnd),
	.combout(\my_reg[17][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[17][12]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[17][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N16
cycloneive_lcell_comb \my_reg[23][12]~feeder (
// Equation(s):
// \my_reg[23][12]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat21),
	.cin(gnd),
	.combout(\my_reg[23][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[23][12]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[23][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N30
cycloneive_lcell_comb \my_reg[9][9]~feeder (
// Equation(s):
// \my_reg[9][9]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat24),
	.cin(gnd),
	.combout(\my_reg[9][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[9][9]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[9][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N28
cycloneive_lcell_comb \my_reg[17][9]~feeder (
// Equation(s):
// \my_reg[17][9]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat24),
	.cin(gnd),
	.combout(\my_reg[17][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[17][9]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[17][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N12
cycloneive_lcell_comb \my_reg[30][9]~feeder (
// Equation(s):
// \my_reg[30][9]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat24),
	.cin(gnd),
	.combout(\my_reg[30][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[30][9]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[30][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N26
cycloneive_lcell_comb \my_reg[21][8]~feeder (
// Equation(s):
// \my_reg[21][8]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat25),
	.cin(gnd),
	.combout(\my_reg[21][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][8]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[21][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N10
cycloneive_lcell_comb \my_reg[22][8]~feeder (
// Equation(s):
// \my_reg[22][8]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat25),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[22][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[22][8]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[22][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N26
cycloneive_lcell_comb \my_reg[24][7]~feeder (
// Equation(s):
// \my_reg[24][7]~feeder_combout  = \wdat~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat26),
	.cin(gnd),
	.combout(\my_reg[24][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[24][7]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[24][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N12
cycloneive_lcell_comb \my_reg[19][7]~feeder (
// Equation(s):
// \my_reg[19][7]~feeder_combout  = \wdat~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat26),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[19][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[19][7]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[19][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N16
cycloneive_lcell_comb \my_reg[1][6]~feeder (
// Equation(s):
// \my_reg[1][6]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat27),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[1][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[1][6]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[1][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N26
cycloneive_lcell_comb \my_reg[17][6]~feeder (
// Equation(s):
// \my_reg[17][6]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat27),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[17][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[17][6]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[17][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N26
cycloneive_lcell_comb \my_reg[25][5]~feeder (
// Equation(s):
// \my_reg[25][5]~feeder_combout  = \wdat~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat28),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[25][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][5]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[25][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N2
cycloneive_lcell_comb \my_reg[26][5]~feeder (
// Equation(s):
// \my_reg[26][5]~feeder_combout  = \wdat~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat28),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[26][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[26][5]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[26][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N6
cycloneive_lcell_comb \my_reg[24][3]~feeder (
// Equation(s):
// \my_reg[24][3]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat30),
	.cin(gnd),
	.combout(\my_reg[24][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[24][3]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[24][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N4
cycloneive_lcell_comb \my_reg[16][3]~feeder (
// Equation(s):
// \my_reg[16][3]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat30),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[16][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[16][3]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[16][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N30
cycloneive_lcell_comb \my_reg[20][2]~feeder (
// Equation(s):
// \my_reg[20][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat31),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[20][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[20][2]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[20][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N20
cycloneive_lcell_comb \my_reg[10][2]~feeder (
// Equation(s):
// \my_reg[10][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat31),
	.cin(gnd),
	.combout(\my_reg[10][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[10][2]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[10][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N0
cycloneive_lcell_comb \Mux63~9 (
// Equation(s):
// Mux63 = (dcifimemload_16 & ((\Mux63~6_combout  & ((\Mux63~8_combout ))) # (!\Mux63~6_combout  & (\Mux63~1_combout )))) # (!dcifimemload_16 & (((\Mux63~6_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux63~1_combout ),
	.datac(\Mux63~6_combout ),
	.datad(\Mux63~8_combout ),
	.cin(gnd),
	.combout(Mux63),
	.cout());
// synopsys translate_off
defparam \Mux63~9 .lut_mask = 16'hF858;
defparam \Mux63~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N14
cycloneive_lcell_comb \Mux63~23 (
// Equation(s):
// Mux631 = (dcifimemload_19 & ((\Mux63~20_combout  & (\Mux63~22_combout )) # (!\Mux63~20_combout  & ((\Mux63~11_combout ))))) # (!dcifimemload_19 & (\Mux63~20_combout ))

	.dataa(dcifimemload_19),
	.datab(\Mux63~20_combout ),
	.datac(\Mux63~22_combout ),
	.datad(\Mux63~11_combout ),
	.cin(gnd),
	.combout(Mux631),
	.cout());
// synopsys translate_off
defparam \Mux63~23 .lut_mask = 16'hE6C4;
defparam \Mux63~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N26
cycloneive_lcell_comb \Mux30~9 (
// Equation(s):
// Mux30 = (dcifimemload_21 & ((\Mux30~6_combout  & ((\Mux30~8_combout ))) # (!\Mux30~6_combout  & (\Mux30~1_combout )))) # (!dcifimemload_21 & (((\Mux30~6_combout ))))

	.dataa(\Mux30~1_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux30~6_combout ),
	.datad(\Mux30~8_combout ),
	.cin(gnd),
	.combout(Mux30),
	.cout());
// synopsys translate_off
defparam \Mux30~9 .lut_mask = 16'hF838;
defparam \Mux30~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N2
cycloneive_lcell_comb \Mux30~19 (
// Equation(s):
// Mux301 = (dcifimemload_24 & ((\Mux30~16_combout  & ((\Mux30~18_combout ))) # (!\Mux30~16_combout  & (\Mux30~11_combout )))) # (!dcifimemload_24 & (\Mux30~16_combout ))

	.dataa(dcifimemload_24),
	.datab(\Mux30~16_combout ),
	.datac(\Mux30~11_combout ),
	.datad(\Mux30~18_combout ),
	.cin(gnd),
	.combout(Mux301),
	.cout());
// synopsys translate_off
defparam \Mux30~19 .lut_mask = 16'hEC64;
defparam \Mux30~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N12
cycloneive_lcell_comb \Mux30~20 (
// Equation(s):
// Mux302 = (dcifimemload_25 & (Mux30)) # (!dcifimemload_25 & ((Mux301)))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(Mux30),
	.datad(Mux301),
	.cin(gnd),
	.combout(Mux302),
	.cout());
// synopsys translate_off
defparam \Mux30~20 .lut_mask = 16'hF3C0;
defparam \Mux30~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N28
cycloneive_lcell_comb \Mux0~20 (
// Equation(s):
// Mux0 = (dcifimemload_25 & (\Mux0~9_combout )) # (!dcifimemload_25 & ((\Mux0~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux0~9_combout ),
	.datad(\Mux0~19_combout ),
	.cin(gnd),
	.combout(Mux0),
	.cout());
// synopsys translate_off
defparam \Mux0~20 .lut_mask = 16'hF5A0;
defparam \Mux0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N10
cycloneive_lcell_comb \Mux32~9 (
// Equation(s):
// Mux32 = (dcifimemload_18 & ((\Mux32~6_combout  & ((\Mux32~8_combout ))) # (!\Mux32~6_combout  & (\Mux32~1_combout )))) # (!dcifimemload_18 & (((\Mux32~6_combout ))))

	.dataa(\Mux32~1_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux32~8_combout ),
	.datad(\Mux32~6_combout ),
	.cin(gnd),
	.combout(Mux32),
	.cout());
// synopsys translate_off
defparam \Mux32~9 .lut_mask = 16'hF388;
defparam \Mux32~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N24
cycloneive_lcell_comb \Mux32~19 (
// Equation(s):
// Mux321 = (dcifimemload_16 & ((\Mux32~16_combout  & (\Mux32~18_combout )) # (!\Mux32~16_combout  & ((\Mux32~11_combout ))))) # (!dcifimemload_16 & (((\Mux32~16_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux32~18_combout ),
	.datac(\Mux32~11_combout ),
	.datad(\Mux32~16_combout ),
	.cin(gnd),
	.combout(Mux321),
	.cout());
// synopsys translate_off
defparam \Mux32~19 .lut_mask = 16'hDDA0;
defparam \Mux32~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N24
cycloneive_lcell_comb \Mux1~20 (
// Equation(s):
// Mux1 = (dcifimemload_25 & (\Mux1~9_combout )) # (!dcifimemload_25 & ((\Mux1~19_combout )))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux1~9_combout ),
	.datad(\Mux1~19_combout ),
	.cin(gnd),
	.combout(Mux1),
	.cout());
// synopsys translate_off
defparam \Mux1~20 .lut_mask = 16'hF3C0;
defparam \Mux1~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N4
cycloneive_lcell_comb \Mux33~9 (
// Equation(s):
// Mux33 = (dcifimemload_19 & ((\Mux33~6_combout  & ((\Mux33~8_combout ))) # (!\Mux33~6_combout  & (\Mux33~1_combout )))) # (!dcifimemload_19 & (((\Mux33~6_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux33~1_combout ),
	.datac(\Mux33~6_combout ),
	.datad(\Mux33~8_combout ),
	.cin(gnd),
	.combout(Mux33),
	.cout());
// synopsys translate_off
defparam \Mux33~9 .lut_mask = 16'hF858;
defparam \Mux33~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N10
cycloneive_lcell_comb \Mux33~19 (
// Equation(s):
// Mux331 = (dcifimemload_16 & ((\Mux33~16_combout  & ((\Mux33~18_combout ))) # (!\Mux33~16_combout  & (\Mux33~11_combout )))) # (!dcifimemload_16 & (((\Mux33~16_combout ))))

	.dataa(\Mux33~11_combout ),
	.datab(\Mux33~18_combout ),
	.datac(dcifimemload_16),
	.datad(\Mux33~16_combout ),
	.cin(gnd),
	.combout(Mux331),
	.cout());
// synopsys translate_off
defparam \Mux33~19 .lut_mask = 16'hCFA0;
defparam \Mux33~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N2
cycloneive_lcell_comb \Mux2~20 (
// Equation(s):
// Mux2 = (dcifimemload_25 & ((\Mux2~9_combout ))) # (!dcifimemload_25 & (\Mux2~19_combout ))

	.dataa(dcifimemload_25),
	.datab(\Mux2~19_combout ),
	.datac(\Mux2~9_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(Mux2),
	.cout());
// synopsys translate_off
defparam \Mux2~20 .lut_mask = 16'hE4E4;
defparam \Mux2~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N20
cycloneive_lcell_comb \Mux34~9 (
// Equation(s):
// Mux34 = (dcifimemload_18 & ((\Mux34~6_combout  & ((\Mux34~8_combout ))) # (!\Mux34~6_combout  & (\Mux34~1_combout )))) # (!dcifimemload_18 & (((\Mux34~6_combout ))))

	.dataa(\Mux34~1_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux34~8_combout ),
	.datad(\Mux34~6_combout ),
	.cin(gnd),
	.combout(Mux34),
	.cout());
// synopsys translate_off
defparam \Mux34~9 .lut_mask = 16'hF388;
defparam \Mux34~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N8
cycloneive_lcell_comb \Mux34~19 (
// Equation(s):
// Mux341 = (dcifimemload_16 & ((\Mux34~16_combout  & ((\Mux34~18_combout ))) # (!\Mux34~16_combout  & (\Mux34~11_combout )))) # (!dcifimemload_16 & (((\Mux34~16_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux34~11_combout ),
	.datac(\Mux34~16_combout ),
	.datad(\Mux34~18_combout ),
	.cin(gnd),
	.combout(Mux341),
	.cout());
// synopsys translate_off
defparam \Mux34~19 .lut_mask = 16'hF858;
defparam \Mux34~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N22
cycloneive_lcell_comb \Mux3~20 (
// Equation(s):
// Mux3 = (dcifimemload_25 & ((\Mux3~9_combout ))) # (!dcifimemload_25 & (\Mux3~19_combout ))

	.dataa(dcifimemload_25),
	.datab(\Mux3~19_combout ),
	.datac(gnd),
	.datad(\Mux3~9_combout ),
	.cin(gnd),
	.combout(Mux3),
	.cout());
// synopsys translate_off
defparam \Mux3~20 .lut_mask = 16'hEE44;
defparam \Mux3~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N6
cycloneive_lcell_comb \Mux35~9 (
// Equation(s):
// Mux35 = (dcifimemload_19 & ((\Mux35~6_combout  & (\Mux35~8_combout )) # (!\Mux35~6_combout  & ((\Mux35~1_combout ))))) # (!dcifimemload_19 & (((\Mux35~6_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux35~8_combout ),
	.datac(\Mux35~6_combout ),
	.datad(\Mux35~1_combout ),
	.cin(gnd),
	.combout(Mux35),
	.cout());
// synopsys translate_off
defparam \Mux35~9 .lut_mask = 16'hDAD0;
defparam \Mux35~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N4
cycloneive_lcell_comb \Mux35~19 (
// Equation(s):
// Mux351 = (\Mux35~16_combout  & (((\Mux35~18_combout ) # (!dcifimemload_16)))) # (!\Mux35~16_combout  & (\Mux35~11_combout  & ((dcifimemload_16))))

	.dataa(\Mux35~11_combout ),
	.datab(\Mux35~18_combout ),
	.datac(\Mux35~16_combout ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(Mux351),
	.cout());
// synopsys translate_off
defparam \Mux35~19 .lut_mask = 16'hCAF0;
defparam \Mux35~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N2
cycloneive_lcell_comb \Mux4~20 (
// Equation(s):
// Mux4 = (dcifimemload_25 & (\Mux4~9_combout )) # (!dcifimemload_25 & ((\Mux4~19_combout )))

	.dataa(\Mux4~9_combout ),
	.datab(dcifimemload_25),
	.datac(gnd),
	.datad(\Mux4~19_combout ),
	.cin(gnd),
	.combout(Mux4),
	.cout());
// synopsys translate_off
defparam \Mux4~20 .lut_mask = 16'hBB88;
defparam \Mux4~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N16
cycloneive_lcell_comb \Mux36~9 (
// Equation(s):
// Mux36 = (dcifimemload_18 & ((\Mux36~6_combout  & (\Mux36~8_combout )) # (!\Mux36~6_combout  & ((\Mux36~1_combout ))))) # (!dcifimemload_18 & (((\Mux36~6_combout ))))

	.dataa(dcifimemload_18),
	.datab(\Mux36~8_combout ),
	.datac(\Mux36~1_combout ),
	.datad(\Mux36~6_combout ),
	.cin(gnd),
	.combout(Mux36),
	.cout());
// synopsys translate_off
defparam \Mux36~9 .lut_mask = 16'hDDA0;
defparam \Mux36~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N6
cycloneive_lcell_comb \Mux36~19 (
// Equation(s):
// Mux361 = (dcifimemload_16 & ((\Mux36~16_combout  & ((\Mux36~18_combout ))) # (!\Mux36~16_combout  & (\Mux36~11_combout )))) # (!dcifimemload_16 & (((\Mux36~16_combout ))))

	.dataa(\Mux36~11_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux36~18_combout ),
	.datad(\Mux36~16_combout ),
	.cin(gnd),
	.combout(Mux361),
	.cout());
// synopsys translate_off
defparam \Mux36~19 .lut_mask = 16'hF388;
defparam \Mux36~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N18
cycloneive_lcell_comb \Mux5~20 (
// Equation(s):
// Mux5 = (dcifimemload_25 & (\Mux5~9_combout )) # (!dcifimemload_25 & ((\Mux5~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux5~9_combout ),
	.datad(\Mux5~19_combout ),
	.cin(gnd),
	.combout(Mux5),
	.cout());
// synopsys translate_off
defparam \Mux5~20 .lut_mask = 16'hF5A0;
defparam \Mux5~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N14
cycloneive_lcell_comb \Mux37~9 (
// Equation(s):
// Mux37 = (dcifimemload_19 & ((\Mux37~6_combout  & (\Mux37~8_combout )) # (!\Mux37~6_combout  & ((\Mux37~1_combout ))))) # (!dcifimemload_19 & (((\Mux37~6_combout ))))

	.dataa(\Mux37~8_combout ),
	.datab(dcifimemload_19),
	.datac(\Mux37~1_combout ),
	.datad(\Mux37~6_combout ),
	.cin(gnd),
	.combout(Mux37),
	.cout());
// synopsys translate_off
defparam \Mux37~9 .lut_mask = 16'hBBC0;
defparam \Mux37~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N8
cycloneive_lcell_comb \Mux37~19 (
// Equation(s):
// Mux371 = (dcifimemload_16 & ((\Mux37~16_combout  & (\Mux37~18_combout )) # (!\Mux37~16_combout  & ((\Mux37~11_combout ))))) # (!dcifimemload_16 & (((\Mux37~16_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux37~18_combout ),
	.datac(\Mux37~11_combout ),
	.datad(\Mux37~16_combout ),
	.cin(gnd),
	.combout(Mux371),
	.cout());
// synopsys translate_off
defparam \Mux37~19 .lut_mask = 16'hDDA0;
defparam \Mux37~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N4
cycloneive_lcell_comb \Mux6~20 (
// Equation(s):
// Mux6 = (dcifimemload_25 & ((\Mux6~9_combout ))) # (!dcifimemload_25 & (\Mux6~19_combout ))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux6~19_combout ),
	.datad(\Mux6~9_combout ),
	.cin(gnd),
	.combout(Mux6),
	.cout());
// synopsys translate_off
defparam \Mux6~20 .lut_mask = 16'hFC30;
defparam \Mux6~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N28
cycloneive_lcell_comb \Mux38~9 (
// Equation(s):
// Mux38 = (\Mux38~6_combout  & (((\Mux38~8_combout )) # (!dcifimemload_18))) # (!\Mux38~6_combout  & (dcifimemload_18 & ((\Mux38~1_combout ))))

	.dataa(\Mux38~6_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux38~8_combout ),
	.datad(\Mux38~1_combout ),
	.cin(gnd),
	.combout(Mux38),
	.cout());
// synopsys translate_off
defparam \Mux38~9 .lut_mask = 16'hE6A2;
defparam \Mux38~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N22
cycloneive_lcell_comb \Mux38~19 (
// Equation(s):
// Mux381 = (dcifimemload_16 & ((\Mux38~16_combout  & ((\Mux38~18_combout ))) # (!\Mux38~16_combout  & (\Mux38~11_combout )))) # (!dcifimemload_16 & (((\Mux38~16_combout ))))

	.dataa(\Mux38~11_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux38~18_combout ),
	.datad(\Mux38~16_combout ),
	.cin(gnd),
	.combout(Mux381),
	.cout());
// synopsys translate_off
defparam \Mux38~19 .lut_mask = 16'hF388;
defparam \Mux38~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N6
cycloneive_lcell_comb \Mux7~9 (
// Equation(s):
// Mux7 = (dcifimemload_21 & ((\Mux7~6_combout  & ((\Mux7~8_combout ))) # (!\Mux7~6_combout  & (\Mux7~1_combout )))) # (!dcifimemload_21 & (((\Mux7~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux7~1_combout ),
	.datac(\Mux7~8_combout ),
	.datad(\Mux7~6_combout ),
	.cin(gnd),
	.combout(Mux7),
	.cout());
// synopsys translate_off
defparam \Mux7~9 .lut_mask = 16'hF588;
defparam \Mux7~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N26
cycloneive_lcell_comb \Mux7~19 (
// Equation(s):
// Mux71 = (dcifimemload_23 & ((\Mux7~16_combout  & ((\Mux7~18_combout ))) # (!\Mux7~16_combout  & (\Mux7~11_combout )))) # (!dcifimemload_23 & (((\Mux7~16_combout ))))

	.dataa(dcifimemload_23),
	.datab(\Mux7~11_combout ),
	.datac(\Mux7~18_combout ),
	.datad(\Mux7~16_combout ),
	.cin(gnd),
	.combout(Mux71),
	.cout());
// synopsys translate_off
defparam \Mux7~19 .lut_mask = 16'hF588;
defparam \Mux7~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N4
cycloneive_lcell_comb \Mux7~20 (
// Equation(s):
// Mux72 = (dcifimemload_25 & ((Mux7))) # (!dcifimemload_25 & (Mux71))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(Mux71),
	.datad(Mux7),
	.cin(gnd),
	.combout(Mux72),
	.cout());
// synopsys translate_off
defparam \Mux7~20 .lut_mask = 16'hFC30;
defparam \Mux7~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N4
cycloneive_lcell_comb \Mux39~9 (
// Equation(s):
// Mux39 = (\Mux39~6_combout  & (((\Mux39~8_combout )) # (!dcifimemload_19))) # (!\Mux39~6_combout  & (dcifimemload_19 & ((\Mux39~1_combout ))))

	.dataa(\Mux39~6_combout ),
	.datab(dcifimemload_19),
	.datac(\Mux39~8_combout ),
	.datad(\Mux39~1_combout ),
	.cin(gnd),
	.combout(Mux39),
	.cout());
// synopsys translate_off
defparam \Mux39~9 .lut_mask = 16'hE6A2;
defparam \Mux39~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N10
cycloneive_lcell_comb \Mux39~19 (
// Equation(s):
// Mux391 = (dcifimemload_16 & ((\Mux39~16_combout  & ((\Mux39~18_combout ))) # (!\Mux39~16_combout  & (\Mux39~11_combout )))) # (!dcifimemload_16 & (((\Mux39~16_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux39~11_combout ),
	.datac(\Mux39~18_combout ),
	.datad(\Mux39~16_combout ),
	.cin(gnd),
	.combout(Mux391),
	.cout());
// synopsys translate_off
defparam \Mux39~19 .lut_mask = 16'hF588;
defparam \Mux39~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N12
cycloneive_lcell_comb \Mux8~20 (
// Equation(s):
// Mux8 = (dcifimemload_25 & ((\Mux8~9_combout ))) # (!dcifimemload_25 & (\Mux8~19_combout ))

	.dataa(dcifimemload_25),
	.datab(\Mux8~19_combout ),
	.datac(gnd),
	.datad(\Mux8~9_combout ),
	.cin(gnd),
	.combout(Mux8),
	.cout());
// synopsys translate_off
defparam \Mux8~20 .lut_mask = 16'hEE44;
defparam \Mux8~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N26
cycloneive_lcell_comb \Mux40~9 (
// Equation(s):
// Mux40 = (dcifimemload_18 & ((\Mux40~6_combout  & ((\Mux40~8_combout ))) # (!\Mux40~6_combout  & (\Mux40~1_combout )))) # (!dcifimemload_18 & (((\Mux40~6_combout ))))

	.dataa(\Mux40~1_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux40~6_combout ),
	.datad(\Mux40~8_combout ),
	.cin(gnd),
	.combout(Mux40),
	.cout());
// synopsys translate_off
defparam \Mux40~9 .lut_mask = 16'hF838;
defparam \Mux40~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N14
cycloneive_lcell_comb \Mux40~19 (
// Equation(s):
// Mux401 = (dcifimemload_16 & ((\Mux40~16_combout  & (\Mux40~18_combout )) # (!\Mux40~16_combout  & ((\Mux40~11_combout ))))) # (!dcifimemload_16 & (((\Mux40~16_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux40~18_combout ),
	.datac(\Mux40~11_combout ),
	.datad(\Mux40~16_combout ),
	.cin(gnd),
	.combout(Mux401),
	.cout());
// synopsys translate_off
defparam \Mux40~19 .lut_mask = 16'hDDA0;
defparam \Mux40~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N2
cycloneive_lcell_comb \Mux9~20 (
// Equation(s):
// Mux9 = (dcifimemload_25 & ((\Mux9~9_combout ))) # (!dcifimemload_25 & (\Mux9~19_combout ))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux9~19_combout ),
	.datad(\Mux9~9_combout ),
	.cin(gnd),
	.combout(Mux9),
	.cout());
// synopsys translate_off
defparam \Mux9~20 .lut_mask = 16'hFA50;
defparam \Mux9~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N22
cycloneive_lcell_comb \Mux41~9 (
// Equation(s):
// Mux41 = (dcifimemload_19 & ((\Mux41~6_combout  & ((\Mux41~8_combout ))) # (!\Mux41~6_combout  & (\Mux41~1_combout )))) # (!dcifimemload_19 & (((\Mux41~6_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux41~1_combout ),
	.datac(\Mux41~6_combout ),
	.datad(\Mux41~8_combout ),
	.cin(gnd),
	.combout(Mux41),
	.cout());
// synopsys translate_off
defparam \Mux41~9 .lut_mask = 16'hF858;
defparam \Mux41~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N16
cycloneive_lcell_comb \Mux41~19 (
// Equation(s):
// Mux411 = (dcifimemload_16 & ((\Mux41~16_combout  & (\Mux41~18_combout )) # (!\Mux41~16_combout  & ((\Mux41~11_combout ))))) # (!dcifimemload_16 & (((\Mux41~16_combout ))))

	.dataa(\Mux41~18_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux41~11_combout ),
	.datad(\Mux41~16_combout ),
	.cin(gnd),
	.combout(Mux411),
	.cout());
// synopsys translate_off
defparam \Mux41~19 .lut_mask = 16'hBBC0;
defparam \Mux41~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N8
cycloneive_lcell_comb \Mux10~20 (
// Equation(s):
// Mux10 = (dcifimemload_25 & ((\Mux10~9_combout ))) # (!dcifimemload_25 & (\Mux10~19_combout ))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux10~19_combout ),
	.datad(\Mux10~9_combout ),
	.cin(gnd),
	.combout(Mux10),
	.cout());
// synopsys translate_off
defparam \Mux10~20 .lut_mask = 16'hFA50;
defparam \Mux10~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N18
cycloneive_lcell_comb \Mux42~9 (
// Equation(s):
// Mux42 = (\Mux42~6_combout  & (((\Mux42~8_combout ) # (!dcifimemload_18)))) # (!\Mux42~6_combout  & (\Mux42~1_combout  & (dcifimemload_18)))

	.dataa(\Mux42~6_combout ),
	.datab(\Mux42~1_combout ),
	.datac(dcifimemload_18),
	.datad(\Mux42~8_combout ),
	.cin(gnd),
	.combout(Mux42),
	.cout());
// synopsys translate_off
defparam \Mux42~9 .lut_mask = 16'hEA4A;
defparam \Mux42~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N8
cycloneive_lcell_comb \Mux42~19 (
// Equation(s):
// Mux421 = (dcifimemload_16 & ((\Mux42~16_combout  & ((\Mux42~18_combout ))) # (!\Mux42~16_combout  & (\Mux42~11_combout )))) # (!dcifimemload_16 & (((\Mux42~16_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux42~11_combout ),
	.datac(\Mux42~16_combout ),
	.datad(\Mux42~18_combout ),
	.cin(gnd),
	.combout(Mux421),
	.cout());
// synopsys translate_off
defparam \Mux42~19 .lut_mask = 16'hF858;
defparam \Mux42~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N20
cycloneive_lcell_comb \Mux11~20 (
// Equation(s):
// Mux11 = (dcifimemload_25 & ((\Mux11~9_combout ))) # (!dcifimemload_25 & (\Mux11~19_combout ))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux11~19_combout ),
	.datad(\Mux11~9_combout ),
	.cin(gnd),
	.combout(Mux11),
	.cout());
// synopsys translate_off
defparam \Mux11~20 .lut_mask = 16'hFA50;
defparam \Mux11~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N8
cycloneive_lcell_comb \Mux43~9 (
// Equation(s):
// Mux43 = (dcifimemload_19 & ((\Mux43~6_combout  & ((\Mux43~8_combout ))) # (!\Mux43~6_combout  & (\Mux43~1_combout )))) # (!dcifimemload_19 & (((\Mux43~6_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux43~1_combout ),
	.datac(\Mux43~6_combout ),
	.datad(\Mux43~8_combout ),
	.cin(gnd),
	.combout(Mux43),
	.cout());
// synopsys translate_off
defparam \Mux43~9 .lut_mask = 16'hF858;
defparam \Mux43~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N16
cycloneive_lcell_comb \Mux43~19 (
// Equation(s):
// Mux431 = (dcifimemload_16 & ((\Mux43~16_combout  & (\Mux43~18_combout )) # (!\Mux43~16_combout  & ((\Mux43~11_combout ))))) # (!dcifimemload_16 & (((\Mux43~16_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux43~18_combout ),
	.datac(\Mux43~11_combout ),
	.datad(\Mux43~16_combout ),
	.cin(gnd),
	.combout(Mux431),
	.cout());
// synopsys translate_off
defparam \Mux43~19 .lut_mask = 16'hDDA0;
defparam \Mux43~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N16
cycloneive_lcell_comb \Mux12~20 (
// Equation(s):
// Mux12 = (dcifimemload_25 & (\Mux12~9_combout )) # (!dcifimemload_25 & ((\Mux12~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux12~9_combout ),
	.datad(\Mux12~19_combout ),
	.cin(gnd),
	.combout(Mux12),
	.cout());
// synopsys translate_off
defparam \Mux12~20 .lut_mask = 16'hF5A0;
defparam \Mux12~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N26
cycloneive_lcell_comb \Mux44~9 (
// Equation(s):
// Mux44 = (\Mux44~6_combout  & (((\Mux44~8_combout )) # (!dcifimemload_18))) # (!\Mux44~6_combout  & (dcifimemload_18 & ((\Mux44~1_combout ))))

	.dataa(\Mux44~6_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux44~8_combout ),
	.datad(\Mux44~1_combout ),
	.cin(gnd),
	.combout(Mux44),
	.cout());
// synopsys translate_off
defparam \Mux44~9 .lut_mask = 16'hE6A2;
defparam \Mux44~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N4
cycloneive_lcell_comb \Mux44~19 (
// Equation(s):
// Mux441 = (dcifimemload_16 & ((\Mux44~16_combout  & ((\Mux44~18_combout ))) # (!\Mux44~16_combout  & (\Mux44~11_combout )))) # (!dcifimemload_16 & (((\Mux44~16_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux44~11_combout ),
	.datac(\Mux44~18_combout ),
	.datad(\Mux44~16_combout ),
	.cin(gnd),
	.combout(Mux441),
	.cout());
// synopsys translate_off
defparam \Mux44~19 .lut_mask = 16'hF588;
defparam \Mux44~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N2
cycloneive_lcell_comb \Mux13~20 (
// Equation(s):
// Mux13 = (dcifimemload_25 & ((\Mux13~9_combout ))) # (!dcifimemload_25 & (\Mux13~19_combout ))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux13~19_combout ),
	.datad(\Mux13~9_combout ),
	.cin(gnd),
	.combout(Mux13),
	.cout());
// synopsys translate_off
defparam \Mux13~20 .lut_mask = 16'hFA50;
defparam \Mux13~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N14
cycloneive_lcell_comb \Mux45~9 (
// Equation(s):
// Mux45 = (dcifimemload_19 & ((\Mux45~6_combout  & (\Mux45~8_combout )) # (!\Mux45~6_combout  & ((\Mux45~1_combout ))))) # (!dcifimemload_19 & (((\Mux45~6_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux45~8_combout ),
	.datac(\Mux45~1_combout ),
	.datad(\Mux45~6_combout ),
	.cin(gnd),
	.combout(Mux45),
	.cout());
// synopsys translate_off
defparam \Mux45~9 .lut_mask = 16'hDDA0;
defparam \Mux45~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N6
cycloneive_lcell_comb \Mux45~19 (
// Equation(s):
// Mux451 = (dcifimemload_16 & ((\Mux45~16_combout  & (\Mux45~18_combout )) # (!\Mux45~16_combout  & ((\Mux45~11_combout ))))) # (!dcifimemload_16 & (((\Mux45~16_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux45~18_combout ),
	.datac(\Mux45~16_combout ),
	.datad(\Mux45~11_combout ),
	.cin(gnd),
	.combout(Mux451),
	.cout());
// synopsys translate_off
defparam \Mux45~19 .lut_mask = 16'hDAD0;
defparam \Mux45~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N0
cycloneive_lcell_comb \Mux14~20 (
// Equation(s):
// Mux14 = (dcifimemload_25 & ((\Mux14~9_combout ))) # (!dcifimemload_25 & (\Mux14~19_combout ))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux14~19_combout ),
	.datad(\Mux14~9_combout ),
	.cin(gnd),
	.combout(Mux14),
	.cout());
// synopsys translate_off
defparam \Mux14~20 .lut_mask = 16'hFA50;
defparam \Mux14~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N24
cycloneive_lcell_comb \Mux46~9 (
// Equation(s):
// Mux46 = (dcifimemload_18 & ((\Mux46~6_combout  & ((\Mux46~8_combout ))) # (!\Mux46~6_combout  & (\Mux46~1_combout )))) # (!dcifimemload_18 & (((\Mux46~6_combout ))))

	.dataa(dcifimemload_18),
	.datab(\Mux46~1_combout ),
	.datac(\Mux46~8_combout ),
	.datad(\Mux46~6_combout ),
	.cin(gnd),
	.combout(Mux46),
	.cout());
// synopsys translate_off
defparam \Mux46~9 .lut_mask = 16'hF588;
defparam \Mux46~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N16
cycloneive_lcell_comb \Mux46~19 (
// Equation(s):
// Mux461 = (dcifimemload_16 & ((\Mux46~16_combout  & ((\Mux46~18_combout ))) # (!\Mux46~16_combout  & (\Mux46~11_combout )))) # (!dcifimemload_16 & (((\Mux46~16_combout ))))

	.dataa(\Mux46~11_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux46~18_combout ),
	.datad(\Mux46~16_combout ),
	.cin(gnd),
	.combout(Mux461),
	.cout());
// synopsys translate_off
defparam \Mux46~19 .lut_mask = 16'hF388;
defparam \Mux46~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N4
cycloneive_lcell_comb \Mux15~20 (
// Equation(s):
// Mux15 = (dcifimemload_25 & ((\Mux15~9_combout ))) # (!dcifimemload_25 & (\Mux15~19_combout ))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux15~19_combout ),
	.datad(\Mux15~9_combout ),
	.cin(gnd),
	.combout(Mux15),
	.cout());
// synopsys translate_off
defparam \Mux15~20 .lut_mask = 16'hFC30;
defparam \Mux15~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N8
cycloneive_lcell_comb \Mux47~9 (
// Equation(s):
// Mux47 = (dcifimemload_19 & ((\Mux47~6_combout  & ((\Mux47~8_combout ))) # (!\Mux47~6_combout  & (\Mux47~1_combout )))) # (!dcifimemload_19 & (((\Mux47~6_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux47~1_combout ),
	.datac(\Mux47~8_combout ),
	.datad(\Mux47~6_combout ),
	.cin(gnd),
	.combout(Mux47),
	.cout());
// synopsys translate_off
defparam \Mux47~9 .lut_mask = 16'hF588;
defparam \Mux47~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N14
cycloneive_lcell_comb \Mux47~19 (
// Equation(s):
// Mux471 = (dcifimemload_16 & ((\Mux47~16_combout  & ((\Mux47~18_combout ))) # (!\Mux47~16_combout  & (\Mux47~11_combout )))) # (!dcifimemload_16 & (((\Mux47~16_combout ))))

	.dataa(\Mux47~11_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux47~16_combout ),
	.datad(\Mux47~18_combout ),
	.cin(gnd),
	.combout(Mux471),
	.cout());
// synopsys translate_off
defparam \Mux47~19 .lut_mask = 16'hF838;
defparam \Mux47~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N16
cycloneive_lcell_comb \Mux16~20 (
// Equation(s):
// Mux16 = (dcifimemload_25 & (\Mux16~9_combout )) # (!dcifimemload_25 & ((\Mux16~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux16~9_combout ),
	.datad(\Mux16~19_combout ),
	.cin(gnd),
	.combout(Mux16),
	.cout());
// synopsys translate_off
defparam \Mux16~20 .lut_mask = 16'hF5A0;
defparam \Mux16~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N16
cycloneive_lcell_comb \Mux48~9 (
// Equation(s):
// Mux48 = (dcifimemload_18 & ((\Mux48~6_combout  & ((\Mux48~8_combout ))) # (!\Mux48~6_combout  & (\Mux48~1_combout )))) # (!dcifimemload_18 & (((\Mux48~6_combout ))))

	.dataa(dcifimemload_18),
	.datab(\Mux48~1_combout ),
	.datac(\Mux48~8_combout ),
	.datad(\Mux48~6_combout ),
	.cin(gnd),
	.combout(Mux48),
	.cout());
// synopsys translate_off
defparam \Mux48~9 .lut_mask = 16'hF588;
defparam \Mux48~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N4
cycloneive_lcell_comb \Mux48~19 (
// Equation(s):
// Mux481 = (dcifimemload_16 & ((\Mux48~16_combout  & (\Mux48~18_combout )) # (!\Mux48~16_combout  & ((\Mux48~11_combout ))))) # (!dcifimemload_16 & (((\Mux48~16_combout ))))

	.dataa(\Mux48~18_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux48~16_combout ),
	.datad(\Mux48~11_combout ),
	.cin(gnd),
	.combout(Mux481),
	.cout());
// synopsys translate_off
defparam \Mux48~19 .lut_mask = 16'hBCB0;
defparam \Mux48~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N6
cycloneive_lcell_comb \Mux17~20 (
// Equation(s):
// Mux17 = (dcifimemload_25 & ((\Mux17~9_combout ))) # (!dcifimemload_25 & (\Mux17~19_combout ))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux17~19_combout ),
	.datad(\Mux17~9_combout ),
	.cin(gnd),
	.combout(Mux17),
	.cout());
// synopsys translate_off
defparam \Mux17~20 .lut_mask = 16'hFA50;
defparam \Mux17~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N0
cycloneive_lcell_comb \Mux49~9 (
// Equation(s):
// Mux49 = (dcifimemload_19 & ((\Mux49~6_combout  & (\Mux49~8_combout )) # (!\Mux49~6_combout  & ((\Mux49~1_combout ))))) # (!dcifimemload_19 & (((\Mux49~6_combout ))))

	.dataa(\Mux49~8_combout ),
	.datab(\Mux49~1_combout ),
	.datac(dcifimemload_19),
	.datad(\Mux49~6_combout ),
	.cin(gnd),
	.combout(Mux49),
	.cout());
// synopsys translate_off
defparam \Mux49~9 .lut_mask = 16'hAFC0;
defparam \Mux49~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N4
cycloneive_lcell_comb \Mux49~19 (
// Equation(s):
// Mux491 = (dcifimemload_16 & ((\Mux49~16_combout  & ((\Mux49~18_combout ))) # (!\Mux49~16_combout  & (\Mux49~11_combout )))) # (!dcifimemload_16 & (((\Mux49~16_combout ))))

	.dataa(\Mux49~11_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux49~16_combout ),
	.datad(\Mux49~18_combout ),
	.cin(gnd),
	.combout(Mux491),
	.cout());
// synopsys translate_off
defparam \Mux49~19 .lut_mask = 16'hF838;
defparam \Mux49~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N0
cycloneive_lcell_comb \Mux18~20 (
// Equation(s):
// Mux18 = (dcifimemload_25 & ((\Mux18~9_combout ))) # (!dcifimemload_25 & (\Mux18~19_combout ))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux18~19_combout ),
	.datad(\Mux18~9_combout ),
	.cin(gnd),
	.combout(Mux18),
	.cout());
// synopsys translate_off
defparam \Mux18~20 .lut_mask = 16'hFC30;
defparam \Mux18~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N16
cycloneive_lcell_comb \Mux50~9 (
// Equation(s):
// Mux50 = (dcifimemload_18 & ((\Mux50~6_combout  & (\Mux50~8_combout )) # (!\Mux50~6_combout  & ((\Mux50~1_combout ))))) # (!dcifimemload_18 & (((\Mux50~6_combout ))))

	.dataa(\Mux50~8_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux50~6_combout ),
	.datad(\Mux50~1_combout ),
	.cin(gnd),
	.combout(Mux50),
	.cout());
// synopsys translate_off
defparam \Mux50~9 .lut_mask = 16'hBCB0;
defparam \Mux50~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N14
cycloneive_lcell_comb \Mux50~19 (
// Equation(s):
// Mux501 = (dcifimemload_16 & ((\Mux50~16_combout  & ((\Mux50~18_combout ))) # (!\Mux50~16_combout  & (\Mux50~11_combout )))) # (!dcifimemload_16 & (((\Mux50~16_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux50~11_combout ),
	.datac(\Mux50~18_combout ),
	.datad(\Mux50~16_combout ),
	.cin(gnd),
	.combout(Mux501),
	.cout());
// synopsys translate_off
defparam \Mux50~19 .lut_mask = 16'hF588;
defparam \Mux50~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N14
cycloneive_lcell_comb \Mux19~20 (
// Equation(s):
// Mux19 = (dcifimemload_25 & (\Mux19~9_combout )) # (!dcifimemload_25 & ((\Mux19~19_combout )))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(\Mux19~9_combout ),
	.datad(\Mux19~19_combout ),
	.cin(gnd),
	.combout(Mux19),
	.cout());
// synopsys translate_off
defparam \Mux19~20 .lut_mask = 16'hF5A0;
defparam \Mux19~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N18
cycloneive_lcell_comb \Mux51~9 (
// Equation(s):
// Mux51 = (dcifimemload_19 & ((\Mux51~6_combout  & ((\Mux51~8_combout ))) # (!\Mux51~6_combout  & (\Mux51~1_combout )))) # (!dcifimemload_19 & (((\Mux51~6_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux51~1_combout ),
	.datac(\Mux51~8_combout ),
	.datad(\Mux51~6_combout ),
	.cin(gnd),
	.combout(Mux51),
	.cout());
// synopsys translate_off
defparam \Mux51~9 .lut_mask = 16'hF588;
defparam \Mux51~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N2
cycloneive_lcell_comb \Mux51~19 (
// Equation(s):
// Mux511 = (dcifimemload_16 & ((\Mux51~16_combout  & ((\Mux51~18_combout ))) # (!\Mux51~16_combout  & (\Mux51~11_combout )))) # (!dcifimemload_16 & (((\Mux51~16_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux51~11_combout ),
	.datac(\Mux51~18_combout ),
	.datad(\Mux51~16_combout ),
	.cin(gnd),
	.combout(Mux511),
	.cout());
// synopsys translate_off
defparam \Mux51~19 .lut_mask = 16'hF588;
defparam \Mux51~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N30
cycloneive_lcell_comb \Mux20~20 (
// Equation(s):
// Mux20 = (dcifimemload_25 & ((\Mux20~9_combout ))) # (!dcifimemload_25 & (\Mux20~19_combout ))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux20~19_combout ),
	.datad(\Mux20~9_combout ),
	.cin(gnd),
	.combout(Mux20),
	.cout());
// synopsys translate_off
defparam \Mux20~20 .lut_mask = 16'hFC30;
defparam \Mux20~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N18
cycloneive_lcell_comb \Mux52~9 (
// Equation(s):
// Mux52 = (dcifimemload_18 & ((\Mux52~6_combout  & (\Mux52~8_combout )) # (!\Mux52~6_combout  & ((\Mux52~1_combout ))))) # (!dcifimemload_18 & (((\Mux52~6_combout ))))

	.dataa(\Mux52~8_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux52~6_combout ),
	.datad(\Mux52~1_combout ),
	.cin(gnd),
	.combout(Mux52),
	.cout());
// synopsys translate_off
defparam \Mux52~9 .lut_mask = 16'hBCB0;
defparam \Mux52~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N0
cycloneive_lcell_comb \Mux52~19 (
// Equation(s):
// Mux521 = (dcifimemload_16 & ((\Mux52~16_combout  & (\Mux52~18_combout )) # (!\Mux52~16_combout  & ((\Mux52~11_combout ))))) # (!dcifimemload_16 & (((\Mux52~16_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux52~18_combout ),
	.datac(\Mux52~11_combout ),
	.datad(\Mux52~16_combout ),
	.cin(gnd),
	.combout(Mux521),
	.cout());
// synopsys translate_off
defparam \Mux52~19 .lut_mask = 16'hDDA0;
defparam \Mux52~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N18
cycloneive_lcell_comb \Mux21~20 (
// Equation(s):
// Mux21 = (dcifimemload_25 & (\Mux21~9_combout )) # (!dcifimemload_25 & ((\Mux21~19_combout )))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux21~9_combout ),
	.datad(\Mux21~19_combout ),
	.cin(gnd),
	.combout(Mux21),
	.cout());
// synopsys translate_off
defparam \Mux21~20 .lut_mask = 16'hF3C0;
defparam \Mux21~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N28
cycloneive_lcell_comb \Mux53~9 (
// Equation(s):
// Mux53 = (dcifimemload_19 & ((\Mux53~6_combout  & ((\Mux53~8_combout ))) # (!\Mux53~6_combout  & (\Mux53~1_combout )))) # (!dcifimemload_19 & (((\Mux53~6_combout ))))

	.dataa(\Mux53~1_combout ),
	.datab(dcifimemload_19),
	.datac(\Mux53~6_combout ),
	.datad(\Mux53~8_combout ),
	.cin(gnd),
	.combout(Mux53),
	.cout());
// synopsys translate_off
defparam \Mux53~9 .lut_mask = 16'hF838;
defparam \Mux53~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N26
cycloneive_lcell_comb \Mux53~19 (
// Equation(s):
// Mux531 = (dcifimemload_16 & ((\Mux53~16_combout  & ((\Mux53~18_combout ))) # (!\Mux53~16_combout  & (\Mux53~11_combout )))) # (!dcifimemload_16 & (((\Mux53~16_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux53~11_combout ),
	.datac(\Mux53~18_combout ),
	.datad(\Mux53~16_combout ),
	.cin(gnd),
	.combout(Mux531),
	.cout());
// synopsys translate_off
defparam \Mux53~19 .lut_mask = 16'hF588;
defparam \Mux53~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N6
cycloneive_lcell_comb \Mux22~20 (
// Equation(s):
// Mux22 = (dcifimemload_25 & (\Mux22~9_combout )) # (!dcifimemload_25 & ((\Mux22~19_combout )))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux22~9_combout ),
	.datad(\Mux22~19_combout ),
	.cin(gnd),
	.combout(Mux22),
	.cout());
// synopsys translate_off
defparam \Mux22~20 .lut_mask = 16'hF3C0;
defparam \Mux22~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N28
cycloneive_lcell_comb \Mux54~9 (
// Equation(s):
// Mux54 = (\Mux54~6_combout  & (((\Mux54~8_combout )) # (!dcifimemload_18))) # (!\Mux54~6_combout  & (dcifimemload_18 & ((\Mux54~1_combout ))))

	.dataa(\Mux54~6_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux54~8_combout ),
	.datad(\Mux54~1_combout ),
	.cin(gnd),
	.combout(Mux54),
	.cout());
// synopsys translate_off
defparam \Mux54~9 .lut_mask = 16'hE6A2;
defparam \Mux54~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N18
cycloneive_lcell_comb \Mux54~19 (
// Equation(s):
// Mux541 = (dcifimemload_16 & ((\Mux54~16_combout  & ((\Mux54~18_combout ))) # (!\Mux54~16_combout  & (\Mux54~11_combout )))) # (!dcifimemload_16 & (((\Mux54~16_combout ))))

	.dataa(\Mux54~11_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux54~18_combout ),
	.datad(\Mux54~16_combout ),
	.cin(gnd),
	.combout(Mux541),
	.cout());
// synopsys translate_off
defparam \Mux54~19 .lut_mask = 16'hF388;
defparam \Mux54~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N14
cycloneive_lcell_comb \Mux23~20 (
// Equation(s):
// Mux23 = (dcifimemload_25 & (\Mux23~9_combout )) # (!dcifimemload_25 & ((\Mux23~19_combout )))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux23~9_combout ),
	.datad(\Mux23~19_combout ),
	.cin(gnd),
	.combout(Mux23),
	.cout());
// synopsys translate_off
defparam \Mux23~20 .lut_mask = 16'hF3C0;
defparam \Mux23~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N0
cycloneive_lcell_comb \Mux55~9 (
// Equation(s):
// Mux55 = (dcifimemload_19 & ((\Mux55~6_combout  & (\Mux55~8_combout )) # (!\Mux55~6_combout  & ((\Mux55~1_combout ))))) # (!dcifimemload_19 & (((\Mux55~6_combout ))))

	.dataa(\Mux55~8_combout ),
	.datab(dcifimemload_19),
	.datac(\Mux55~6_combout ),
	.datad(\Mux55~1_combout ),
	.cin(gnd),
	.combout(Mux55),
	.cout());
// synopsys translate_off
defparam \Mux55~9 .lut_mask = 16'hBCB0;
defparam \Mux55~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N6
cycloneive_lcell_comb \Mux55~19 (
// Equation(s):
// Mux551 = (dcifimemload_16 & ((\Mux55~16_combout  & (\Mux55~18_combout )) # (!\Mux55~16_combout  & ((\Mux55~11_combout ))))) # (!dcifimemload_16 & (((\Mux55~16_combout ))))

	.dataa(\Mux55~18_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux55~16_combout ),
	.datad(\Mux55~11_combout ),
	.cin(gnd),
	.combout(Mux551),
	.cout());
// synopsys translate_off
defparam \Mux55~19 .lut_mask = 16'hBCB0;
defparam \Mux55~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N30
cycloneive_lcell_comb \Mux24~9 (
// Equation(s):
// Mux24 = (dcifimemload_21 & ((\Mux24~6_combout  & (\Mux24~8_combout )) # (!\Mux24~6_combout  & ((\Mux24~1_combout ))))) # (!dcifimemload_21 & (((\Mux24~6_combout ))))

	.dataa(\Mux24~8_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux24~1_combout ),
	.datad(\Mux24~6_combout ),
	.cin(gnd),
	.combout(Mux24),
	.cout());
// synopsys translate_off
defparam \Mux24~9 .lut_mask = 16'hBBC0;
defparam \Mux24~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N24
cycloneive_lcell_comb \Mux24~19 (
// Equation(s):
// Mux241 = (dcifimemload_24 & ((\Mux24~16_combout  & ((\Mux24~18_combout ))) # (!\Mux24~16_combout  & (\Mux24~11_combout )))) # (!dcifimemload_24 & (((\Mux24~16_combout ))))

	.dataa(\Mux24~11_combout ),
	.datab(dcifimemload_24),
	.datac(\Mux24~16_combout ),
	.datad(\Mux24~18_combout ),
	.cin(gnd),
	.combout(Mux241),
	.cout());
// synopsys translate_off
defparam \Mux24~19 .lut_mask = 16'hF838;
defparam \Mux24~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N18
cycloneive_lcell_comb \Mux24~20 (
// Equation(s):
// Mux242 = (dcifimemload_25 & (Mux24)) # (!dcifimemload_25 & ((Mux241)))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(Mux24),
	.datad(Mux241),
	.cin(gnd),
	.combout(Mux242),
	.cout());
// synopsys translate_off
defparam \Mux24~20 .lut_mask = 16'hF3C0;
defparam \Mux24~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N28
cycloneive_lcell_comb \Mux56~9 (
// Equation(s):
// Mux56 = (dcifimemload_18 & ((\Mux56~6_combout  & (\Mux56~8_combout )) # (!\Mux56~6_combout  & ((\Mux56~1_combout ))))) # (!dcifimemload_18 & (((\Mux56~6_combout ))))

	.dataa(dcifimemload_18),
	.datab(\Mux56~8_combout ),
	.datac(\Mux56~6_combout ),
	.datad(\Mux56~1_combout ),
	.cin(gnd),
	.combout(Mux56),
	.cout());
// synopsys translate_off
defparam \Mux56~9 .lut_mask = 16'hDAD0;
defparam \Mux56~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N22
cycloneive_lcell_comb \Mux56~19 (
// Equation(s):
// Mux561 = (dcifimemload_16 & ((\Mux56~16_combout  & (\Mux56~18_combout )) # (!\Mux56~16_combout  & ((\Mux56~11_combout ))))) # (!dcifimemload_16 & (((\Mux56~16_combout ))))

	.dataa(\Mux56~18_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux56~11_combout ),
	.datad(\Mux56~16_combout ),
	.cin(gnd),
	.combout(Mux561),
	.cout());
// synopsys translate_off
defparam \Mux56~19 .lut_mask = 16'hBBC0;
defparam \Mux56~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N16
cycloneive_lcell_comb \Mux25~9 (
// Equation(s):
// Mux25 = (dcifimemload_21 & ((\Mux25~6_combout  & ((\Mux25~8_combout ))) # (!\Mux25~6_combout  & (\Mux25~1_combout )))) # (!dcifimemload_21 & (((\Mux25~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux25~1_combout ),
	.datac(\Mux25~6_combout ),
	.datad(\Mux25~8_combout ),
	.cin(gnd),
	.combout(Mux25),
	.cout());
// synopsys translate_off
defparam \Mux25~9 .lut_mask = 16'hF858;
defparam \Mux25~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N4
cycloneive_lcell_comb \Mux25~19 (
// Equation(s):
// Mux251 = (dcifimemload_23 & ((\Mux25~16_combout  & (\Mux25~18_combout )) # (!\Mux25~16_combout  & ((\Mux25~11_combout ))))) # (!dcifimemload_23 & (((\Mux25~16_combout ))))

	.dataa(\Mux25~18_combout ),
	.datab(dcifimemload_23),
	.datac(\Mux25~11_combout ),
	.datad(\Mux25~16_combout ),
	.cin(gnd),
	.combout(Mux251),
	.cout());
// synopsys translate_off
defparam \Mux25~19 .lut_mask = 16'hBBC0;
defparam \Mux25~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N30
cycloneive_lcell_comb \Mux25~20 (
// Equation(s):
// Mux252 = (dcifimemload_25 & ((Mux25))) # (!dcifimemload_25 & (Mux251))

	.dataa(dcifimemload_25),
	.datab(gnd),
	.datac(Mux251),
	.datad(Mux25),
	.cin(gnd),
	.combout(Mux252),
	.cout());
// synopsys translate_off
defparam \Mux25~20 .lut_mask = 16'hFA50;
defparam \Mux25~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N20
cycloneive_lcell_comb \Mux57~9 (
// Equation(s):
// Mux57 = (dcifimemload_19 & ((\Mux57~6_combout  & ((\Mux57~8_combout ))) # (!\Mux57~6_combout  & (\Mux57~1_combout )))) # (!dcifimemload_19 & (((\Mux57~6_combout ))))

	.dataa(\Mux57~1_combout ),
	.datab(dcifimemload_19),
	.datac(\Mux57~6_combout ),
	.datad(\Mux57~8_combout ),
	.cin(gnd),
	.combout(Mux57),
	.cout());
// synopsys translate_off
defparam \Mux57~9 .lut_mask = 16'hF838;
defparam \Mux57~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N22
cycloneive_lcell_comb \Mux57~19 (
// Equation(s):
// Mux571 = (dcifimemload_16 & ((\Mux57~16_combout  & ((\Mux57~18_combout ))) # (!\Mux57~16_combout  & (\Mux57~11_combout )))) # (!dcifimemload_16 & (((\Mux57~16_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux57~11_combout ),
	.datac(\Mux57~16_combout ),
	.datad(\Mux57~18_combout ),
	.cin(gnd),
	.combout(Mux571),
	.cout());
// synopsys translate_off
defparam \Mux57~19 .lut_mask = 16'hF858;
defparam \Mux57~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N18
cycloneive_lcell_comb \Mux26~20 (
// Equation(s):
// Mux26 = (dcifimemload_25 & ((\Mux26~9_combout ))) # (!dcifimemload_25 & (\Mux26~19_combout ))

	.dataa(\Mux26~19_combout ),
	.datab(dcifimemload_25),
	.datac(gnd),
	.datad(\Mux26~9_combout ),
	.cin(gnd),
	.combout(Mux26),
	.cout());
// synopsys translate_off
defparam \Mux26~20 .lut_mask = 16'hEE22;
defparam \Mux26~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N6
cycloneive_lcell_comb \Mux58~9 (
// Equation(s):
// Mux58 = (dcifimemload_18 & ((\Mux58~6_combout  & ((\Mux58~8_combout ))) # (!\Mux58~6_combout  & (\Mux58~1_combout )))) # (!dcifimemload_18 & (((\Mux58~6_combout ))))

	.dataa(dcifimemload_18),
	.datab(\Mux58~1_combout ),
	.datac(\Mux58~8_combout ),
	.datad(\Mux58~6_combout ),
	.cin(gnd),
	.combout(Mux58),
	.cout());
// synopsys translate_off
defparam \Mux58~9 .lut_mask = 16'hF588;
defparam \Mux58~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N8
cycloneive_lcell_comb \Mux58~19 (
// Equation(s):
// Mux581 = (dcifimemload_16 & ((\Mux58~16_combout  & (\Mux58~18_combout )) # (!\Mux58~16_combout  & ((\Mux58~11_combout ))))) # (!dcifimemload_16 & (((\Mux58~16_combout ))))

	.dataa(\Mux58~18_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux58~16_combout ),
	.datad(\Mux58~11_combout ),
	.cin(gnd),
	.combout(Mux581),
	.cout());
// synopsys translate_off
defparam \Mux58~19 .lut_mask = 16'hBCB0;
defparam \Mux58~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N6
cycloneive_lcell_comb \Mux27~9 (
// Equation(s):
// Mux27 = (dcifimemload_21 & ((\Mux27~6_combout  & ((\Mux27~8_combout ))) # (!\Mux27~6_combout  & (\Mux27~1_combout )))) # (!dcifimemload_21 & (((\Mux27~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux27~1_combout ),
	.datac(\Mux27~8_combout ),
	.datad(\Mux27~6_combout ),
	.cin(gnd),
	.combout(Mux27),
	.cout());
// synopsys translate_off
defparam \Mux27~9 .lut_mask = 16'hF588;
defparam \Mux27~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N0
cycloneive_lcell_comb \Mux27~19 (
// Equation(s):
// Mux271 = (\Mux27~16_combout  & (((\Mux27~18_combout )) # (!dcifimemload_23))) # (!\Mux27~16_combout  & (dcifimemload_23 & ((\Mux27~11_combout ))))

	.dataa(\Mux27~16_combout ),
	.datab(dcifimemload_23),
	.datac(\Mux27~18_combout ),
	.datad(\Mux27~11_combout ),
	.cin(gnd),
	.combout(Mux271),
	.cout());
// synopsys translate_off
defparam \Mux27~19 .lut_mask = 16'hE6A2;
defparam \Mux27~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N26
cycloneive_lcell_comb \Mux27~20 (
// Equation(s):
// Mux272 = (dcifimemload_25 & ((Mux27))) # (!dcifimemload_25 & (Mux271))

	.dataa(gnd),
	.datab(Mux271),
	.datac(dcifimemload_25),
	.datad(Mux27),
	.cin(gnd),
	.combout(Mux272),
	.cout());
// synopsys translate_off
defparam \Mux27~20 .lut_mask = 16'hFC0C;
defparam \Mux27~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N10
cycloneive_lcell_comb \Mux59~9 (
// Equation(s):
// Mux59 = (dcifimemload_19 & ((\Mux59~6_combout  & ((\Mux59~8_combout ))) # (!\Mux59~6_combout  & (\Mux59~1_combout )))) # (!dcifimemload_19 & (((\Mux59~6_combout ))))

	.dataa(\Mux59~1_combout ),
	.datab(\Mux59~8_combout ),
	.datac(dcifimemload_19),
	.datad(\Mux59~6_combout ),
	.cin(gnd),
	.combout(Mux59),
	.cout());
// synopsys translate_off
defparam \Mux59~9 .lut_mask = 16'hCFA0;
defparam \Mux59~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N4
cycloneive_lcell_comb \Mux59~19 (
// Equation(s):
// Mux591 = (dcifimemload_16 & ((\Mux59~16_combout  & (\Mux59~18_combout )) # (!\Mux59~16_combout  & ((\Mux59~11_combout ))))) # (!dcifimemload_16 & (((\Mux59~16_combout ))))

	.dataa(\Mux59~18_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux59~16_combout ),
	.datad(\Mux59~11_combout ),
	.cin(gnd),
	.combout(Mux591),
	.cout());
// synopsys translate_off
defparam \Mux59~19 .lut_mask = 16'hBCB0;
defparam \Mux59~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N0
cycloneive_lcell_comb \Mux28~20 (
// Equation(s):
// Mux28 = (dcifimemload_25 & ((\Mux28~9_combout ))) # (!dcifimemload_25 & (\Mux28~19_combout ))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(\Mux28~19_combout ),
	.datad(\Mux28~9_combout ),
	.cin(gnd),
	.combout(Mux28),
	.cout());
// synopsys translate_off
defparam \Mux28~20 .lut_mask = 16'hFC30;
defparam \Mux28~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N10
cycloneive_lcell_comb \Mux60~9 (
// Equation(s):
// Mux60 = (dcifimemload_16 & ((\Mux60~6_combout  & (\Mux60~8_combout )) # (!\Mux60~6_combout  & ((\Mux60~1_combout ))))) # (!dcifimemload_16 & (((\Mux60~6_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux60~8_combout ),
	.datac(\Mux60~1_combout ),
	.datad(\Mux60~6_combout ),
	.cin(gnd),
	.combout(Mux60),
	.cout());
// synopsys translate_off
defparam \Mux60~9 .lut_mask = 16'hDDA0;
defparam \Mux60~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N30
cycloneive_lcell_comb \Mux60~19 (
// Equation(s):
// Mux601 = (dcifimemload_18 & ((\Mux60~16_combout  & ((\Mux60~18_combout ))) # (!\Mux60~16_combout  & (\Mux60~11_combout )))) # (!dcifimemload_18 & (((\Mux60~16_combout ))))

	.dataa(\Mux60~11_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux60~18_combout ),
	.datad(\Mux60~16_combout ),
	.cin(gnd),
	.combout(Mux601),
	.cout());
// synopsys translate_off
defparam \Mux60~19 .lut_mask = 16'hF388;
defparam \Mux60~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N6
cycloneive_lcell_comb \Mux29~9 (
// Equation(s):
// Mux29 = (dcifimemload_21 & ((\Mux29~6_combout  & (\Mux29~8_combout )) # (!\Mux29~6_combout  & ((\Mux29~1_combout ))))) # (!dcifimemload_21 & (((\Mux29~6_combout ))))

	.dataa(\Mux29~8_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux29~1_combout ),
	.datad(\Mux29~6_combout ),
	.cin(gnd),
	.combout(Mux29),
	.cout());
// synopsys translate_off
defparam \Mux29~9 .lut_mask = 16'hBBC0;
defparam \Mux29~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N4
cycloneive_lcell_comb \Mux29~19 (
// Equation(s):
// Mux291 = (dcifimemload_23 & ((\Mux29~16_combout  & (\Mux29~18_combout )) # (!\Mux29~16_combout  & ((\Mux29~11_combout ))))) # (!dcifimemload_23 & (((\Mux29~16_combout ))))

	.dataa(\Mux29~18_combout ),
	.datab(dcifimemload_23),
	.datac(\Mux29~11_combout ),
	.datad(\Mux29~16_combout ),
	.cin(gnd),
	.combout(Mux291),
	.cout());
// synopsys translate_off
defparam \Mux29~19 .lut_mask = 16'hBBC0;
defparam \Mux29~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N10
cycloneive_lcell_comb \Mux29~20 (
// Equation(s):
// Mux292 = (dcifimemload_25 & ((Mux29))) # (!dcifimemload_25 & (Mux291))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(Mux291),
	.datad(Mux29),
	.cin(gnd),
	.combout(Mux292),
	.cout());
// synopsys translate_off
defparam \Mux29~20 .lut_mask = 16'hFC30;
defparam \Mux29~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N16
cycloneive_lcell_comb \Mux61~9 (
// Equation(s):
// Mux61 = (dcifimemload_19 & ((\Mux61~6_combout  & ((\Mux61~8_combout ))) # (!\Mux61~6_combout  & (\Mux61~1_combout )))) # (!dcifimemload_19 & (((\Mux61~6_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux61~1_combout ),
	.datac(\Mux61~8_combout ),
	.datad(\Mux61~6_combout ),
	.cin(gnd),
	.combout(Mux61),
	.cout());
// synopsys translate_off
defparam \Mux61~9 .lut_mask = 16'hF588;
defparam \Mux61~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N22
cycloneive_lcell_comb \Mux61~19 (
// Equation(s):
// Mux611 = (dcifimemload_16 & ((\Mux61~16_combout  & ((\Mux61~18_combout ))) # (!\Mux61~16_combout  & (\Mux61~11_combout )))) # (!dcifimemload_16 & (((\Mux61~16_combout ))))

	.dataa(\Mux61~11_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux61~18_combout ),
	.datad(\Mux61~16_combout ),
	.cin(gnd),
	.combout(Mux611),
	.cout());
// synopsys translate_off
defparam \Mux61~19 .lut_mask = 16'hF388;
defparam \Mux61~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N22
cycloneive_lcell_comb \Mux62~9 (
// Equation(s):
// Mux62 = (dcifimemload_16 & ((\Mux62~6_combout  & ((\Mux62~8_combout ))) # (!\Mux62~6_combout  & (\Mux62~1_combout )))) # (!dcifimemload_16 & (((\Mux62~6_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux62~1_combout ),
	.datac(\Mux62~8_combout ),
	.datad(\Mux62~6_combout ),
	.cin(gnd),
	.combout(Mux62),
	.cout());
// synopsys translate_off
defparam \Mux62~9 .lut_mask = 16'hF588;
defparam \Mux62~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N10
cycloneive_lcell_comb \Mux62~21 (
// Equation(s):
// Mux621 = (dcifimemload_18 & ((\Mux62~18_combout  & ((\Mux62~20_combout ))) # (!\Mux62~18_combout  & (\Mux62~11_combout )))) # (!dcifimemload_18 & (((\Mux62~18_combout ))))

	.dataa(\Mux62~11_combout ),
	.datab(dcifimemload_18),
	.datac(\Mux62~20_combout ),
	.datad(\Mux62~18_combout ),
	.cin(gnd),
	.combout(Mux621),
	.cout());
// synopsys translate_off
defparam \Mux62~21 .lut_mask = 16'hF388;
defparam \Mux62~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N2
cycloneive_lcell_comb \Mux31~9 (
// Equation(s):
// Mux31 = (dcifimemload_21 & ((\Mux31~6_combout  & ((\Mux31~8_combout ))) # (!\Mux31~6_combout  & (\Mux31~1_combout )))) # (!dcifimemload_21 & (\Mux31~6_combout ))

	.dataa(dcifimemload_21),
	.datab(\Mux31~6_combout ),
	.datac(\Mux31~1_combout ),
	.datad(\Mux31~8_combout ),
	.cin(gnd),
	.combout(Mux31),
	.cout());
// synopsys translate_off
defparam \Mux31~9 .lut_mask = 16'hEC64;
defparam \Mux31~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N30
cycloneive_lcell_comb \Mux31~19 (
// Equation(s):
// Mux311 = (dcifimemload_23 & ((\Mux31~16_combout  & (\Mux31~18_combout )) # (!\Mux31~16_combout  & ((\Mux31~11_combout ))))) # (!dcifimemload_23 & (((\Mux31~16_combout ))))

	.dataa(dcifimemload_23),
	.datab(\Mux31~18_combout ),
	.datac(\Mux31~16_combout ),
	.datad(\Mux31~11_combout ),
	.cin(gnd),
	.combout(Mux311),
	.cout());
// synopsys translate_off
defparam \Mux31~19 .lut_mask = 16'hDAD0;
defparam \Mux31~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N4
cycloneive_lcell_comb \Mux31~20 (
// Equation(s):
// Mux312 = (dcifimemload_25 & ((Mux31))) # (!dcifimemload_25 & (Mux311))

	.dataa(gnd),
	.datab(dcifimemload_25),
	.datac(Mux311),
	.datad(Mux31),
	.cin(gnd),
	.combout(Mux312),
	.cout());
// synopsys translate_off
defparam \Mux31~20 .lut_mask = 16'hFC30;
defparam \Mux31~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N16
cycloneive_lcell_comb \Decoder0~15 (
// Equation(s):
// \Decoder0~15_combout  = (cuifRegWEN1 & (\wsel~1_combout  & \wsel~0_combout ))

	.dataa(cuifRegWEN),
	.datab(gnd),
	.datac(wsel1),
	.datad(wsel),
	.cin(gnd),
	.combout(\Decoder0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~15 .lut_mask = 16'hA000;
defparam \Decoder0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N26
cycloneive_lcell_comb \Decoder0~16 (
// Equation(s):
// \Decoder0~16_combout  = (\wsel~3_combout  & (\wsel~2_combout  & (!\wsel~4_combout  & \Decoder0~15_combout )))

	.dataa(wsel3),
	.datab(wsel2),
	.datac(wsel4),
	.datad(\Decoder0~15_combout ),
	.cin(gnd),
	.combout(\Decoder0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~16 .lut_mask = 16'h0800;
defparam \Decoder0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N5
dffeas \my_reg[29][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][0] .is_wysiwyg = "true";
defparam \my_reg[29][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N8
cycloneive_lcell_comb \my_reg[25][0]~feeder (
// Equation(s):
// \my_reg[25][0]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat),
	.cin(gnd),
	.combout(\my_reg[25][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][0]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[25][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N30
cycloneive_lcell_comb \Decoder0~10 (
// Equation(s):
// \Decoder0~10_combout  = (!\wsel~4_combout  & (\wsel~2_combout  & !\wsel~3_combout ))

	.dataa(wsel4),
	.datab(wsel2),
	.datac(wsel3),
	.datad(gnd),
	.cin(gnd),
	.combout(\Decoder0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~10 .lut_mask = 16'h0404;
defparam \Decoder0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N4
cycloneive_lcell_comb \Decoder0~11 (
// Equation(s):
// \Decoder0~11_combout  = (\wsel~0_combout  & (\wsel~1_combout  & (\Decoder0~10_combout  & cuifRegWEN1)))

	.dataa(wsel),
	.datab(wsel1),
	.datac(\Decoder0~10_combout ),
	.datad(cuifRegWEN),
	.cin(gnd),
	.combout(\Decoder0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~11 .lut_mask = 16'h8000;
defparam \Decoder0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N9
dffeas \my_reg[25][0] (
	.clk(CLK),
	.d(\my_reg[25][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][0] .is_wysiwyg = "true";
defparam \my_reg[25][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N16
cycloneive_lcell_comb \my_reg[21][0]~feeder (
// Equation(s):
// \my_reg[21][0]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[21][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][0]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[21][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N16
cycloneive_lcell_comb \Decoder0~12 (
// Equation(s):
// \Decoder0~12_combout  = (cuifRegWEN1 & (!\wsel~1_combout  & \wsel~0_combout ))

	.dataa(cuifRegWEN),
	.datab(gnd),
	.datac(wsel1),
	.datad(wsel),
	.cin(gnd),
	.combout(\Decoder0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~12 .lut_mask = 16'h0A00;
defparam \Decoder0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N22
cycloneive_lcell_comb \Decoder0~13 (
// Equation(s):
// \Decoder0~13_combout  = (!\wsel~4_combout  & (\wsel~2_combout  & (\wsel~3_combout  & \Decoder0~12_combout )))

	.dataa(wsel4),
	.datab(wsel2),
	.datac(wsel3),
	.datad(\Decoder0~12_combout ),
	.cin(gnd),
	.combout(\Decoder0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~13 .lut_mask = 16'h4000;
defparam \Decoder0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N17
dffeas \my_reg[21][0] (
	.clk(CLK),
	.d(\my_reg[21][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][0] .is_wysiwyg = "true";
defparam \my_reg[21][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N10
cycloneive_lcell_comb \Mux63~0 (
// Equation(s):
// \Mux63~0_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[21][0]~q ))) # (!dcifimemload_18 & (\my_reg[17][0]~q ))))

	.dataa(\my_reg[17][0]~q ),
	.datab(\my_reg[21][0]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux63~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~0 .lut_mask = 16'hFC0A;
defparam \Mux63~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N30
cycloneive_lcell_comb \Mux63~1 (
// Equation(s):
// \Mux63~1_combout  = (dcifimemload_19 & ((\Mux63~0_combout  & (\my_reg[29][0]~q )) # (!\Mux63~0_combout  & ((\my_reg[25][0]~q ))))) # (!dcifimemload_19 & (((\Mux63~0_combout ))))

	.dataa(\my_reg[29][0]~q ),
	.datab(\my_reg[25][0]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux63~0_combout ),
	.cin(gnd),
	.combout(\Mux63~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~1 .lut_mask = 16'hAFC0;
defparam \Mux63~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N6
cycloneive_lcell_comb \Decoder0~19 (
// Equation(s):
// \Decoder0~19_combout  = (\wsel~0_combout  & (cuifRegWEN1 & (\wsel~1_combout  & !\wsel~2_combout )))

	.dataa(wsel),
	.datab(cuifRegWEN),
	.datac(wsel1),
	.datad(wsel2),
	.cin(gnd),
	.combout(\Decoder0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~19 .lut_mask = 16'h0080;
defparam \Decoder0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N10
cycloneive_lcell_comb \Decoder0~22 (
// Equation(s):
// \Decoder0~22_combout  = (\wsel~3_combout  & (\wsel~4_combout  & \Decoder0~19_combout ))

	.dataa(wsel3),
	.datab(gnd),
	.datac(wsel4),
	.datad(\Decoder0~19_combout ),
	.cin(gnd),
	.combout(\Decoder0~22_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~22 .lut_mask = 16'hA000;
defparam \Decoder0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N19
dffeas \my_reg[30][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][0] .is_wysiwyg = "true";
defparam \my_reg[30][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N30
cycloneive_lcell_comb \Decoder0~17 (
// Equation(s):
// \Decoder0~17_combout  = (\wsel~0_combout  & (cuifRegWEN1 & (!\wsel~2_combout  & !\wsel~1_combout )))

	.dataa(wsel),
	.datab(cuifRegWEN),
	.datac(wsel2),
	.datad(wsel1),
	.cin(gnd),
	.combout(\Decoder0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~17 .lut_mask = 16'h0008;
defparam \Decoder0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N6
cycloneive_lcell_comb \Decoder0~21 (
// Equation(s):
// \Decoder0~21_combout  = (\wsel~4_combout  & (!\wsel~3_combout  & \Decoder0~17_combout ))

	.dataa(wsel4),
	.datab(wsel3),
	.datac(gnd),
	.datad(\Decoder0~17_combout ),
	.cin(gnd),
	.combout(\Decoder0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~21 .lut_mask = 16'h2200;
defparam \Decoder0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N25
dffeas \my_reg[18][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][0] .is_wysiwyg = "true";
defparam \my_reg[18][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N8
cycloneive_lcell_comb \Decoder0~20 (
// Equation(s):
// \Decoder0~20_combout  = (!\wsel~3_combout  & (\wsel~4_combout  & \Decoder0~19_combout ))

	.dataa(wsel3),
	.datab(gnd),
	.datac(wsel4),
	.datad(\Decoder0~19_combout ),
	.cin(gnd),
	.combout(\Decoder0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~20 .lut_mask = 16'h5000;
defparam \Decoder0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N3
dffeas \my_reg[26][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][0] .is_wysiwyg = "true";
defparam \my_reg[26][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N2
cycloneive_lcell_comb \Mux63~2 (
// Equation(s):
// \Mux63~2_combout  = (dcifimemload_19 & (((\my_reg[26][0]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[18][0]~q  & ((!dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[18][0]~q ),
	.datac(\my_reg[26][0]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux63~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~2 .lut_mask = 16'hAAE4;
defparam \Mux63~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N8
cycloneive_lcell_comb \Mux63~3 (
// Equation(s):
// \Mux63~3_combout  = (dcifimemload_18 & ((\Mux63~2_combout  & ((\my_reg[30][0]~q ))) # (!\Mux63~2_combout  & (\my_reg[22][0]~q )))) # (!dcifimemload_18 & (((\Mux63~2_combout ))))

	.dataa(\my_reg[22][0]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[30][0]~q ),
	.datad(\Mux63~2_combout ),
	.cin(gnd),
	.combout(\Mux63~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~3 .lut_mask = 16'hF388;
defparam \Mux63~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N30
cycloneive_lcell_comb \Decoder0~24 (
// Equation(s):
// \Decoder0~24_combout  = (!\wsel~4_combout  & (\Decoder0~17_combout  & !\wsel~3_combout ))

	.dataa(gnd),
	.datab(wsel4),
	.datac(\Decoder0~17_combout ),
	.datad(wsel3),
	.cin(gnd),
	.combout(\Decoder0~24_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~24 .lut_mask = 16'h0030;
defparam \Decoder0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N3
dffeas \my_reg[16][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][0] .is_wysiwyg = "true";
defparam \my_reg[16][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N20
cycloneive_lcell_comb \Decoder0~23 (
// Equation(s):
// \Decoder0~23_combout  = (\wsel~3_combout  & (!\wsel~4_combout  & \Decoder0~17_combout ))

	.dataa(wsel3),
	.datab(gnd),
	.datac(wsel4),
	.datad(\Decoder0~17_combout ),
	.cin(gnd),
	.combout(\Decoder0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~23 .lut_mask = 16'h0A00;
defparam \Decoder0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N9
dffeas \my_reg[20][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][0] .is_wysiwyg = "true";
defparam \my_reg[20][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N24
cycloneive_lcell_comb \Decoder0~26 (
// Equation(s):
// \Decoder0~26_combout  = (!\wsel~3_combout  & (!\wsel~4_combout  & \Decoder0~19_combout ))

	.dataa(wsel3),
	.datab(gnd),
	.datac(wsel4),
	.datad(\Decoder0~19_combout ),
	.cin(gnd),
	.combout(\Decoder0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~26 .lut_mask = 16'h0500;
defparam \Decoder0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N19
dffeas \my_reg[24][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][0] .is_wysiwyg = "true";
defparam \my_reg[24][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N18
cycloneive_lcell_comb \Mux63~4 (
// Equation(s):
// \Mux63~4_combout  = (dcifimemload_19 & ((dcifimemload_18 & (\my_reg[28][0]~q )) # (!dcifimemload_18 & ((\my_reg[24][0]~q ))))) # (!dcifimemload_19 & (((dcifimemload_18))))

	.dataa(\my_reg[28][0]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[24][0]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux63~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~4 .lut_mask = 16'hBBC0;
defparam \Mux63~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N8
cycloneive_lcell_comb \Mux63~5 (
// Equation(s):
// \Mux63~5_combout  = (dcifimemload_19 & (((\Mux63~4_combout )))) # (!dcifimemload_19 & ((\Mux63~4_combout  & ((\my_reg[20][0]~q ))) # (!\Mux63~4_combout  & (\my_reg[16][0]~q ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[16][0]~q ),
	.datac(\my_reg[20][0]~q ),
	.datad(\Mux63~4_combout ),
	.cin(gnd),
	.combout(\Mux63~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~5 .lut_mask = 16'hFA44;
defparam \Mux63~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N26
cycloneive_lcell_comb \Mux63~6 (
// Equation(s):
// \Mux63~6_combout  = (dcifimemload_17 & ((\Mux63~3_combout ) # ((dcifimemload_16)))) # (!dcifimemload_17 & (((!dcifimemload_16 & \Mux63~5_combout ))))

	.dataa(dcifimemload_17),
	.datab(\Mux63~3_combout ),
	.datac(dcifimemload_16),
	.datad(\Mux63~5_combout ),
	.cin(gnd),
	.combout(\Mux63~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~6 .lut_mask = 16'hADA8;
defparam \Mux63~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N20
cycloneive_lcell_comb \Decoder0~30 (
// Equation(s):
// \Decoder0~30_combout  = (\wsel~2_combout  & (\wsel~3_combout  & (\wsel~4_combout  & \Decoder0~15_combout )))

	.dataa(wsel2),
	.datab(wsel3),
	.datac(wsel4),
	.datad(\Decoder0~15_combout ),
	.cin(gnd),
	.combout(\Decoder0~30_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~30 .lut_mask = 16'h8000;
defparam \Decoder0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N21
dffeas \my_reg[31][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][0] .is_wysiwyg = "true";
defparam \my_reg[31][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N28
cycloneive_lcell_comb \my_reg[27][0]~feeder (
// Equation(s):
// \my_reg[27][0]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat),
	.cin(gnd),
	.combout(\my_reg[27][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[27][0]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[27][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N18
cycloneive_lcell_comb \Decoder0~27 (
// Equation(s):
// \Decoder0~27_combout  = (!\wsel~3_combout  & (\wsel~2_combout  & (\wsel~4_combout  & \Decoder0~15_combout )))

	.dataa(wsel3),
	.datab(wsel2),
	.datac(wsel4),
	.datad(\Decoder0~15_combout ),
	.cin(gnd),
	.combout(\Decoder0~27_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~27 .lut_mask = 16'h4000;
defparam \Decoder0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y34_N29
dffeas \my_reg[27][0] (
	.clk(CLK),
	.d(\my_reg[27][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][0] .is_wysiwyg = "true";
defparam \my_reg[27][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N16
cycloneive_lcell_comb \my_reg[23][0]~feeder (
// Equation(s):
// \my_reg[23][0]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[23][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[23][0]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[23][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N28
cycloneive_lcell_comb \Decoder0~28 (
// Equation(s):
// \Decoder0~28_combout  = (\wsel~4_combout  & (\wsel~2_combout  & (\wsel~3_combout  & \Decoder0~12_combout )))

	.dataa(wsel4),
	.datab(wsel2),
	.datac(wsel3),
	.datad(\Decoder0~12_combout ),
	.cin(gnd),
	.combout(\Decoder0~28_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~28 .lut_mask = 16'h8000;
defparam \Decoder0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N17
dffeas \my_reg[23][0] (
	.clk(CLK),
	.d(\my_reg[23][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][0] .is_wysiwyg = "true";
defparam \my_reg[23][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N18
cycloneive_lcell_comb \Mux63~7 (
// Equation(s):
// \Mux63~7_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[23][0]~q ))) # (!dcifimemload_18 & (\my_reg[19][0]~q ))))

	.dataa(\my_reg[19][0]~q ),
	.datab(\my_reg[23][0]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux63~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~7 .lut_mask = 16'hFC0A;
defparam \Mux63~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N20
cycloneive_lcell_comb \Mux63~8 (
// Equation(s):
// \Mux63~8_combout  = (dcifimemload_19 & ((\Mux63~7_combout  & (\my_reg[31][0]~q )) # (!\Mux63~7_combout  & ((\my_reg[27][0]~q ))))) # (!dcifimemload_19 & (((\Mux63~7_combout ))))

	.dataa(\my_reg[31][0]~q ),
	.datab(\my_reg[27][0]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux63~7_combout ),
	.cin(gnd),
	.combout(\Mux63~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~8 .lut_mask = 16'hAFC0;
defparam \Mux63~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N10
cycloneive_lcell_comb \Decoder0~51 (
// Equation(s):
// \Decoder0~51_combout  = (\wsel~4_combout  & (!\wsel~0_combout  & (!\wsel~1_combout  & cuifRegWEN1)))

	.dataa(wsel4),
	.datab(wsel),
	.datac(wsel1),
	.datad(cuifRegWEN),
	.cin(gnd),
	.combout(\Decoder0~51_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~51 .lut_mask = 16'h0200;
defparam \Decoder0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N2
cycloneive_lcell_comb \Decoder0~42 (
// Equation(s):
// \Decoder0~42_combout  = (!\wsel~2_combout  & (!\wsel~3_combout  & \Decoder0~51_combout ))

	.dataa(gnd),
	.datab(wsel2),
	.datac(wsel3),
	.datad(\Decoder0~51_combout ),
	.cin(gnd),
	.combout(\Decoder0~42_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~42 .lut_mask = 16'h0300;
defparam \Decoder0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y37_N31
dffeas \my_reg[2][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][0] .is_wysiwyg = "true";
defparam \my_reg[2][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N0
cycloneive_lcell_comb \Decoder0~41 (
// Equation(s):
// \Decoder0~41_combout  = (\wsel~2_combout  & (!\wsel~3_combout  & \Decoder0~51_combout ))

	.dataa(gnd),
	.datab(wsel2),
	.datac(wsel3),
	.datad(\Decoder0~51_combout ),
	.cin(gnd),
	.combout(\Decoder0~41_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~41 .lut_mask = 16'h0C00;
defparam \Decoder0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y37_N1
dffeas \my_reg[3][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][0] .is_wysiwyg = "true";
defparam \my_reg[3][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N20
cycloneive_lcell_comb \Decoder0~52 (
// Equation(s):
// \Decoder0~52_combout  = (!\wsel~0_combout  & (!\wsel~1_combout  & (cuifRegWEN1 & \Decoder0~10_combout )))

	.dataa(wsel),
	.datab(wsel1),
	.datac(cuifRegWEN),
	.datad(\Decoder0~10_combout ),
	.cin(gnd),
	.combout(\Decoder0~52_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~52 .lut_mask = 16'h1000;
defparam \Decoder0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N19
dffeas \my_reg[1][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][0] .is_wysiwyg = "true";
defparam \my_reg[1][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N18
cycloneive_lcell_comb \Mux63~17 (
// Equation(s):
// \Mux63~17_combout  = (ramiframload_17 & (\my_reg[3][0]~q )) # (!ramiframload_17 & ((\my_reg[1][0]~q )))

	.dataa(gnd),
	.datab(\my_reg[3][0]~q ),
	.datac(\my_reg[1][0]~q ),
	.datad(ramiframload_17),
	.cin(gnd),
	.combout(\Mux63~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~17 .lut_mask = 16'hCCF0;
defparam \Mux63~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N4
cycloneive_lcell_comb \Mux63~18 (
// Equation(s):
// \Mux63~18_combout  = (ccifiwait_0 & (((\Mux63~17_combout  & ramiframload_16)))) # (!ccifiwait_0 & (\Mux63~16_combout ))

	.dataa(\Mux63~16_combout ),
	.datab(\Mux63~17_combout ),
	.datac(ccifiwait_0),
	.datad(ramiframload_16),
	.cin(gnd),
	.combout(\Mux63~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~18 .lut_mask = 16'hCA0A;
defparam \Mux63~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N26
cycloneive_lcell_comb \Mux63~19 (
// Equation(s):
// \Mux63~19_combout  = (\Mux63~18_combout ) # ((dcifimemload_17 & (\my_reg[2][0]~q  & !dcifimemload_16)))

	.dataa(dcifimemload_17),
	.datab(\my_reg[2][0]~q ),
	.datac(\Mux63~18_combout ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux63~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~19 .lut_mask = 16'hF0F8;
defparam \Mux63~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N12
cycloneive_lcell_comb \Decoder0~36 (
// Equation(s):
// \Decoder0~36_combout  = (!\wsel~2_combout  & (\wsel~3_combout  & \Decoder0~51_combout ))

	.dataa(gnd),
	.datab(wsel2),
	.datac(wsel3),
	.datad(\Decoder0~51_combout ),
	.cin(gnd),
	.combout(\Decoder0~36_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~36 .lut_mask = 16'h3000;
defparam \Decoder0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N17
dffeas \my_reg[6][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][0] .is_wysiwyg = "true";
defparam \my_reg[6][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N26
cycloneive_lcell_comb \Decoder0~40 (
// Equation(s):
// \Decoder0~40_combout  = (\wsel~2_combout  & (\wsel~3_combout  & \Decoder0~51_combout ))

	.dataa(gnd),
	.datab(wsel2),
	.datac(wsel3),
	.datad(\Decoder0~51_combout ),
	.cin(gnd),
	.combout(\Decoder0~40_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~40 .lut_mask = 16'hC000;
defparam \Decoder0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N17
dffeas \my_reg[7][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][0] .is_wysiwyg = "true";
defparam \my_reg[7][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N16
cycloneive_lcell_comb \Decoder0~35 (
// Equation(s):
// \Decoder0~35_combout  = (!\wsel~1_combout  & !\wsel~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(wsel1),
	.datad(wsel),
	.cin(gnd),
	.combout(\Decoder0~35_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~35 .lut_mask = 16'h000F;
defparam \Decoder0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N6
cycloneive_lcell_comb \Decoder0~37 (
// Equation(s):
// \Decoder0~37_combout  = (cuifRegWEN1 & (!\wsel~4_combout  & (\wsel~3_combout  & \Decoder0~35_combout )))

	.dataa(cuifRegWEN),
	.datab(wsel4),
	.datac(wsel3),
	.datad(\Decoder0~35_combout ),
	.cin(gnd),
	.combout(\Decoder0~37_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~37 .lut_mask = 16'h2000;
defparam \Decoder0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N18
cycloneive_lcell_comb \Decoder0~38 (
// Equation(s):
// \Decoder0~38_combout  = (\wsel~2_combout  & \Decoder0~37_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(wsel2),
	.datad(\Decoder0~37_combout ),
	.cin(gnd),
	.combout(\Decoder0~38_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~38 .lut_mask = 16'hF000;
defparam \Decoder0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N15
dffeas \my_reg[5][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][0] .is_wysiwyg = "true";
defparam \my_reg[5][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N18
cycloneive_lcell_comb \Mux63~13 (
// Equation(s):
// \Mux63~13_combout  = (ramiframload_17 & (((ramiframload_16)))) # (!ramiframload_17 & ((ramiframload_16 & ((\my_reg[5][0]~q ))) # (!ramiframload_16 & (\my_reg[4][0]~q ))))

	.dataa(\my_reg[4][0]~q ),
	.datab(ramiframload_17),
	.datac(\my_reg[5][0]~q ),
	.datad(ramiframload_16),
	.cin(gnd),
	.combout(\Mux63~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~13 .lut_mask = 16'hFC22;
defparam \Mux63~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N6
cycloneive_lcell_comb \Mux63~14 (
// Equation(s):
// \Mux63~14_combout  = (ccifiwait_0 & ((\Mux63~13_combout ))) # (!ccifiwait_0 & (\Mux63~12_combout ))

	.dataa(\Mux63~12_combout ),
	.datab(gnd),
	.datac(ccifiwait_0),
	.datad(\Mux63~13_combout ),
	.cin(gnd),
	.combout(\Mux63~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~14 .lut_mask = 16'hFA0A;
defparam \Mux63~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N16
cycloneive_lcell_comb \Mux63~15 (
// Equation(s):
// \Mux63~15_combout  = (dcifimemload_17 & ((\Mux63~14_combout  & ((\my_reg[7][0]~q ))) # (!\Mux63~14_combout  & (\my_reg[6][0]~q )))) # (!dcifimemload_17 & (((\Mux63~14_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[6][0]~q ),
	.datac(\my_reg[7][0]~q ),
	.datad(\Mux63~14_combout ),
	.cin(gnd),
	.combout(\Mux63~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~15 .lut_mask = 16'hF588;
defparam \Mux63~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N24
cycloneive_lcell_comb \Mux63~20 (
// Equation(s):
// \Mux63~20_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & ((\Mux63~15_combout ))) # (!dcifimemload_18 & (\Mux63~19_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux63~19_combout ),
	.datad(\Mux63~15_combout ),
	.cin(gnd),
	.combout(\Mux63~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~20 .lut_mask = 16'hDC98;
defparam \Mux63~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N20
cycloneive_lcell_comb \my_reg[14][0]~feeder (
// Equation(s):
// \my_reg[14][0]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[14][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[14][0]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[14][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N4
cycloneive_lcell_comb \Decoder0~49 (
// Equation(s):
// \Decoder0~49_combout  = (\wsel~1_combout  & (\wsel~4_combout  & (!\wsel~0_combout  & cuifRegWEN1)))

	.dataa(wsel1),
	.datab(wsel4),
	.datac(wsel),
	.datad(cuifRegWEN),
	.cin(gnd),
	.combout(\Decoder0~49_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~49 .lut_mask = 16'h0800;
defparam \Decoder0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N8
cycloneive_lcell_comb \Decoder0~43 (
// Equation(s):
// \Decoder0~43_combout  = (!\wsel~2_combout  & (\Decoder0~49_combout  & \wsel~3_combout ))

	.dataa(wsel2),
	.datab(gnd),
	.datac(\Decoder0~49_combout ),
	.datad(wsel3),
	.cin(gnd),
	.combout(\Decoder0~43_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~43 .lut_mask = 16'h5000;
defparam \Decoder0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N21
dffeas \my_reg[14][0] (
	.clk(CLK),
	.d(\my_reg[14][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][0] .is_wysiwyg = "true";
defparam \my_reg[14][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N26
cycloneive_lcell_comb \Decoder0~47 (
// Equation(s):
// \Decoder0~47_combout  = (\wsel~2_combout  & (\Decoder0~49_combout  & \wsel~3_combout ))

	.dataa(wsel2),
	.datab(gnd),
	.datac(\Decoder0~49_combout ),
	.datad(wsel3),
	.cin(gnd),
	.combout(\Decoder0~47_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~47 .lut_mask = 16'hA000;
defparam \Decoder0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N1
dffeas \my_reg[15][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][0] .is_wysiwyg = "true";
defparam \my_reg[15][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N8
cycloneive_lcell_comb \my_reg[12][0]~feeder (
// Equation(s):
// \my_reg[12][0]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[12][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[12][0]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[12][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N10
cycloneive_lcell_comb \Decoder0~31 (
// Equation(s):
// \Decoder0~31_combout  = (\wsel~1_combout  & !\wsel~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(wsel1),
	.datad(wsel),
	.cin(gnd),
	.combout(\Decoder0~31_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~31 .lut_mask = 16'h00F0;
defparam \Decoder0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N4
cycloneive_lcell_comb \Decoder0~44 (
// Equation(s):
// \Decoder0~44_combout  = (cuifRegWEN1 & (!\wsel~4_combout  & (\Decoder0~31_combout  & \wsel~3_combout )))

	.dataa(cuifRegWEN),
	.datab(wsel4),
	.datac(\Decoder0~31_combout ),
	.datad(wsel3),
	.cin(gnd),
	.combout(\Decoder0~44_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~44 .lut_mask = 16'h2000;
defparam \Decoder0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N26
cycloneive_lcell_comb \Decoder0~46 (
// Equation(s):
// \Decoder0~46_combout  = (\Decoder0~44_combout  & !\wsel~2_combout )

	.dataa(gnd),
	.datab(\Decoder0~44_combout ),
	.datac(gnd),
	.datad(wsel2),
	.cin(gnd),
	.combout(\Decoder0~46_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~46 .lut_mask = 16'h00CC;
defparam \Decoder0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N9
dffeas \my_reg[12][0] (
	.clk(CLK),
	.d(\my_reg[12][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][0] .is_wysiwyg = "true";
defparam \my_reg[12][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N18
cycloneive_lcell_comb \Decoder0~45 (
// Equation(s):
// \Decoder0~45_combout  = (\Decoder0~44_combout  & \wsel~2_combout )

	.dataa(gnd),
	.datab(\Decoder0~44_combout ),
	.datac(gnd),
	.datad(wsel2),
	.cin(gnd),
	.combout(\Decoder0~45_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~45 .lut_mask = 16'hCC00;
defparam \Decoder0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N5
dffeas \my_reg[13][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][0] .is_wysiwyg = "true";
defparam \my_reg[13][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N2
cycloneive_lcell_comb \Mux63~21 (
// Equation(s):
// \Mux63~21_combout  = (dcifimemload_16 & (((dcifimemload_17) # (\my_reg[13][0]~q )))) # (!dcifimemload_16 & (\my_reg[12][0]~q  & (!dcifimemload_17)))

	.dataa(dcifimemload_16),
	.datab(\my_reg[12][0]~q ),
	.datac(dcifimemload_17),
	.datad(\my_reg[13][0]~q ),
	.cin(gnd),
	.combout(\Mux63~21_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~21 .lut_mask = 16'hAEA4;
defparam \Mux63~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N0
cycloneive_lcell_comb \Mux63~22 (
// Equation(s):
// \Mux63~22_combout  = (dcifimemload_17 & ((\Mux63~21_combout  & ((\my_reg[15][0]~q ))) # (!\Mux63~21_combout  & (\my_reg[14][0]~q )))) # (!dcifimemload_17 & (((\Mux63~21_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[14][0]~q ),
	.datac(\my_reg[15][0]~q ),
	.datad(\Mux63~21_combout ),
	.cin(gnd),
	.combout(\Mux63~22_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~22 .lut_mask = 16'hF588;
defparam \Mux63~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N14
cycloneive_lcell_comb \Decoder0~34 (
// Equation(s):
// \Decoder0~34_combout  = (\wsel~2_combout  & (\Decoder0~49_combout  & !\wsel~3_combout ))

	.dataa(wsel2),
	.datab(gnd),
	.datac(\Decoder0~49_combout ),
	.datad(wsel3),
	.cin(gnd),
	.combout(\Decoder0~34_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~34 .lut_mask = 16'h00A0;
defparam \Decoder0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N15
dffeas \my_reg[11][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][0] .is_wysiwyg = "true";
defparam \my_reg[11][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N22
cycloneive_lcell_comb \my_reg[10][0]~feeder (
// Equation(s):
// \my_reg[10][0]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[10][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[10][0]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[10][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N6
cycloneive_lcell_comb \Decoder0~32 (
// Equation(s):
// \Decoder0~32_combout  = (!\wsel~2_combout  & (\Decoder0~49_combout  & !\wsel~3_combout ))

	.dataa(wsel2),
	.datab(gnd),
	.datac(\Decoder0~49_combout ),
	.datad(wsel3),
	.cin(gnd),
	.combout(\Decoder0~32_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~32 .lut_mask = 16'h0050;
defparam \Decoder0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y42_N23
dffeas \my_reg[10][0] (
	.clk(CLK),
	.d(\my_reg[10][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][0] .is_wysiwyg = "true";
defparam \my_reg[10][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N16
cycloneive_lcell_comb \Mux63~10 (
// Equation(s):
// \Mux63~10_combout  = (dcifimemload_17 & (((\my_reg[10][0]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\my_reg[8][0]~q  & ((!dcifimemload_16))))

	.dataa(\my_reg[8][0]~q ),
	.datab(\my_reg[10][0]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux63~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~10 .lut_mask = 16'hF0CA;
defparam \Mux63~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N4
cycloneive_lcell_comb \Decoder0~48 (
// Equation(s):
// \Decoder0~48_combout  = (cuifRegWEN1 & (\wsel~1_combout  & (\Decoder0~10_combout  & !\wsel~0_combout )))

	.dataa(cuifRegWEN),
	.datab(wsel1),
	.datac(\Decoder0~10_combout ),
	.datad(wsel),
	.cin(gnd),
	.combout(\Decoder0~48_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~48 .lut_mask = 16'h0080;
defparam \Decoder0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y42_N5
dffeas \my_reg[9][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][0] .is_wysiwyg = "true";
defparam \my_reg[9][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N4
cycloneive_lcell_comb \Mux63~11 (
// Equation(s):
// \Mux63~11_combout  = (\Mux63~10_combout  & ((\my_reg[11][0]~q ) # ((!dcifimemload_16)))) # (!\Mux63~10_combout  & (((\my_reg[9][0]~q  & dcifimemload_16))))

	.dataa(\my_reg[11][0]~q ),
	.datab(\Mux63~10_combout ),
	.datac(\my_reg[9][0]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux63~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~11 .lut_mask = 16'hB8CC;
defparam \Mux63~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N17
dffeas \my_reg[25][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][1] .is_wysiwyg = "true";
defparam \my_reg[25][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N8
cycloneive_lcell_comb \my_reg[29][1]~feeder (
// Equation(s):
// \my_reg[29][1]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\my_reg[29][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[29][1]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[29][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N9
dffeas \my_reg[29][1] (
	.clk(CLK),
	.d(\my_reg[29][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][1] .is_wysiwyg = "true";
defparam \my_reg[29][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N31
dffeas \my_reg[21][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][1] .is_wysiwyg = "true";
defparam \my_reg[21][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N16
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\my_reg[21][1]~q ))) # (!dcifimemload_23 & (\my_reg[17][1]~q ))))

	.dataa(\my_reg[17][1]~q ),
	.datab(\my_reg[21][1]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'hFC0A;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N6
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// \Mux30~1_combout  = (dcifimemload_24 & ((\Mux30~0_combout  & ((\my_reg[29][1]~q ))) # (!\Mux30~0_combout  & (\my_reg[25][1]~q )))) # (!dcifimemload_24 & (((\Mux30~0_combout ))))

	.dataa(\my_reg[25][1]~q ),
	.datab(\my_reg[29][1]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux30~0_combout ),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'hCFA0;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N4
cycloneive_lcell_comb \my_reg[20][1]~feeder (
// Equation(s):
// \my_reg[20][1]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\my_reg[20][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[20][1]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[20][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y29_N5
dffeas \my_reg[20][1] (
	.clk(CLK),
	.d(\my_reg[20][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][1] .is_wysiwyg = "true";
defparam \my_reg[20][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N31
dffeas \my_reg[16][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][1] .is_wysiwyg = "true";
defparam \my_reg[16][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N30
cycloneive_lcell_comb \Mux30~4 (
// Equation(s):
// \Mux30~4_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[24][1]~q )) # (!dcifimemload_24 & ((\my_reg[16][1]~q )))))

	.dataa(\my_reg[24][1]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[16][1]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux30~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~4 .lut_mask = 16'hEE30;
defparam \Mux30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N22
cycloneive_lcell_comb \Mux30~5 (
// Equation(s):
// \Mux30~5_combout  = (dcifimemload_23 & ((\Mux30~4_combout  & (\my_reg[28][1]~q )) # (!\Mux30~4_combout  & ((\my_reg[20][1]~q ))))) # (!dcifimemload_23 & (((\Mux30~4_combout ))))

	.dataa(\my_reg[28][1]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[20][1]~q ),
	.datad(\Mux30~4_combout ),
	.cin(gnd),
	.combout(\Mux30~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~5 .lut_mask = 16'hBBC0;
defparam \Mux30~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N5
dffeas \my_reg[30][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][1] .is_wysiwyg = "true";
defparam \my_reg[30][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N17
dffeas \my_reg[18][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][1] .is_wysiwyg = "true";
defparam \my_reg[18][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N16
cycloneive_lcell_comb \Mux30~2 (
// Equation(s):
// \Mux30~2_combout  = (dcifimemload_24 & ((\my_reg[26][1]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\my_reg[18][1]~q  & !dcifimemload_23))))

	.dataa(\my_reg[26][1]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[18][1]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~2 .lut_mask = 16'hCCB8;
defparam \Mux30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N2
cycloneive_lcell_comb \Mux30~3 (
// Equation(s):
// \Mux30~3_combout  = (dcifimemload_23 & ((\Mux30~2_combout  & ((\my_reg[30][1]~q ))) # (!\Mux30~2_combout  & (\my_reg[22][1]~q )))) # (!dcifimemload_23 & (((\Mux30~2_combout ))))

	.dataa(\my_reg[22][1]~q ),
	.datab(\my_reg[30][1]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux30~2_combout ),
	.cin(gnd),
	.combout(\Mux30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~3 .lut_mask = 16'hCFA0;
defparam \Mux30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N4
cycloneive_lcell_comb \Mux30~6 (
// Equation(s):
// \Mux30~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux30~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & (\Mux30~5_combout )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux30~5_combout ),
	.datad(\Mux30~3_combout ),
	.cin(gnd),
	.combout(\Mux30~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~6 .lut_mask = 16'hBA98;
defparam \Mux30~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N26
cycloneive_lcell_comb \my_reg[27][1]~feeder (
// Equation(s):
// \my_reg[27][1]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\my_reg[27][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[27][1]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[27][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y34_N27
dffeas \my_reg[27][1] (
	.clk(CLK),
	.d(\my_reg[27][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][1] .is_wysiwyg = "true";
defparam \my_reg[27][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N3
dffeas \my_reg[31][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][1] .is_wysiwyg = "true";
defparam \my_reg[31][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N25
dffeas \my_reg[23][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][1] .is_wysiwyg = "true";
defparam \my_reg[23][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N24
cycloneive_lcell_comb \Mux30~7 (
// Equation(s):
// \Mux30~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\my_reg[23][1]~q ))) # (!dcifimemload_23 & (\my_reg[19][1]~q ))))

	.dataa(\my_reg[19][1]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[23][1]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux30~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~7 .lut_mask = 16'hFC22;
defparam \Mux30~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N10
cycloneive_lcell_comb \Mux30~8 (
// Equation(s):
// \Mux30~8_combout  = (dcifimemload_24 & ((\Mux30~7_combout  & ((\my_reg[31][1]~q ))) # (!\Mux30~7_combout  & (\my_reg[27][1]~q )))) # (!dcifimemload_24 & (((\Mux30~7_combout ))))

	.dataa(\my_reg[27][1]~q ),
	.datab(\my_reg[31][1]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux30~7_combout ),
	.cin(gnd),
	.combout(\Mux30~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~8 .lut_mask = 16'hCFA0;
defparam \Mux30~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y32_N27
dffeas \my_reg[3][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][1] .is_wysiwyg = "true";
defparam \my_reg[3][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N16
cycloneive_lcell_comb \my_reg[1][1]~feeder (
// Equation(s):
// \my_reg[1][1]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat1),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[1][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[1][1]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[1][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N17
dffeas \my_reg[1][1] (
	.clk(CLK),
	.d(\my_reg[1][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][1] .is_wysiwyg = "true";
defparam \my_reg[1][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N28
cycloneive_lcell_comb \Mux30~14 (
// Equation(s):
// \Mux30~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\my_reg[3][1]~q )) # (!dcifimemload_22 & ((\my_reg[1][1]~q )))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[3][1]~q ),
	.datac(\my_reg[1][1]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux30~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~14 .lut_mask = 16'hD800;
defparam \Mux30~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N15
dffeas \my_reg[2][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][1] .is_wysiwyg = "true";
defparam \my_reg[2][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N14
cycloneive_lcell_comb \Mux30~15 (
// Equation(s):
// \Mux30~15_combout  = (\Mux30~14_combout ) # ((dcifimemload_22 & (\my_reg[2][1]~q  & !dcifimemload_21)))

	.dataa(dcifimemload_22),
	.datab(\Mux30~14_combout ),
	.datac(\my_reg[2][1]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux30~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~15 .lut_mask = 16'hCCEC;
defparam \Mux30~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N13
dffeas \my_reg[6][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][1] .is_wysiwyg = "true";
defparam \my_reg[6][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N27
dffeas \my_reg[7][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][1] .is_wysiwyg = "true";
defparam \my_reg[7][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N7
dffeas \my_reg[5][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][1] .is_wysiwyg = "true";
defparam \my_reg[5][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N28
cycloneive_lcell_comb \Decoder0~39 (
// Equation(s):
// \Decoder0~39_combout  = (!\wsel~2_combout  & \Decoder0~37_combout )

	.dataa(gnd),
	.datab(wsel2),
	.datac(gnd),
	.datad(\Decoder0~37_combout ),
	.cin(gnd),
	.combout(\Decoder0~39_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~39 .lut_mask = 16'h3300;
defparam \Decoder0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N13
dffeas \my_reg[4][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][1] .is_wysiwyg = "true";
defparam \my_reg[4][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N12
cycloneive_lcell_comb \Mux30~12 (
// Equation(s):
// \Mux30~12_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\my_reg[5][1]~q )) # (!dcifimemload_21 & ((\my_reg[4][1]~q )))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[5][1]~q ),
	.datac(\my_reg[4][1]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux30~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~12 .lut_mask = 16'hEE50;
defparam \Mux30~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N26
cycloneive_lcell_comb \Mux30~13 (
// Equation(s):
// \Mux30~13_combout  = (dcifimemload_22 & ((\Mux30~12_combout  & ((\my_reg[7][1]~q ))) # (!\Mux30~12_combout  & (\my_reg[6][1]~q )))) # (!dcifimemload_22 & (((\Mux30~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[6][1]~q ),
	.datac(\my_reg[7][1]~q ),
	.datad(\Mux30~12_combout ),
	.cin(gnd),
	.combout(\Mux30~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~13 .lut_mask = 16'hF588;
defparam \Mux30~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N24
cycloneive_lcell_comb \Mux30~16 (
// Equation(s):
// \Mux30~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & ((\Mux30~13_combout ))) # (!dcifimemload_23 & (\Mux30~15_combout ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux30~15_combout ),
	.datad(\Mux30~13_combout ),
	.cin(gnd),
	.combout(\Mux30~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~16 .lut_mask = 16'hDC98;
defparam \Mux30~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N4
cycloneive_lcell_comb \my_reg[9][1]~feeder (
// Equation(s):
// \my_reg[9][1]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat1),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[9][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[9][1]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[9][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N5
dffeas \my_reg[9][1] (
	.clk(CLK),
	.d(\my_reg[9][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][1] .is_wysiwyg = "true";
defparam \my_reg[9][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N11
dffeas \my_reg[11][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][1] .is_wysiwyg = "true";
defparam \my_reg[11][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N0
cycloneive_lcell_comb \my_reg[10][1]~feeder (
// Equation(s):
// \my_reg[10][1]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\my_reg[10][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[10][1]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[10][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N1
dffeas \my_reg[10][1] (
	.clk(CLK),
	.d(\my_reg[10][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][1] .is_wysiwyg = "true";
defparam \my_reg[10][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N20
cycloneive_lcell_comb \Decoder0~33 (
// Equation(s):
// \Decoder0~33_combout  = (\Decoder0~50_combout  & (!\wsel~4_combout  & (!\wsel~2_combout  & !\wsel~3_combout )))

	.dataa(\Decoder0~50_combout ),
	.datab(wsel4),
	.datac(wsel2),
	.datad(wsel3),
	.cin(gnd),
	.combout(\Decoder0~33_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~33 .lut_mask = 16'h0002;
defparam \Decoder0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N17
dffeas \my_reg[8][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][1] .is_wysiwyg = "true";
defparam \my_reg[8][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N6
cycloneive_lcell_comb \Mux30~10 (
// Equation(s):
// \Mux30~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][1]~q )) # (!dcifimemload_22 & ((\my_reg[8][1]~q )))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[10][1]~q ),
	.datac(\my_reg[8][1]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux30~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~10 .lut_mask = 16'hEE50;
defparam \Mux30~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N20
cycloneive_lcell_comb \Mux30~11 (
// Equation(s):
// \Mux30~11_combout  = (dcifimemload_21 & ((\Mux30~10_combout  & ((\my_reg[11][1]~q ))) # (!\Mux30~10_combout  & (\my_reg[9][1]~q )))) # (!dcifimemload_21 & (((\Mux30~10_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][1]~q ),
	.datac(\my_reg[11][1]~q ),
	.datad(\Mux30~10_combout ),
	.cin(gnd),
	.combout(\Mux30~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~11 .lut_mask = 16'hF588;
defparam \Mux30~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N7
dffeas \my_reg[15][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][1] .is_wysiwyg = "true";
defparam \my_reg[15][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y41_N1
dffeas \my_reg[14][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][1] .is_wysiwyg = "true";
defparam \my_reg[14][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N20
cycloneive_lcell_comb \my_reg[13][1]~feeder (
// Equation(s):
// \my_reg[13][1]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\my_reg[13][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[13][1]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[13][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N21
dffeas \my_reg[13][1] (
	.clk(CLK),
	.d(\my_reg[13][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][1] .is_wysiwyg = "true";
defparam \my_reg[13][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N14
cycloneive_lcell_comb \Mux30~17 (
// Equation(s):
// \Mux30~17_combout  = (dcifimemload_21 & (((\my_reg[13][1]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\my_reg[12][1]~q  & ((!dcifimemload_22))))

	.dataa(\my_reg[12][1]~q ),
	.datab(\my_reg[13][1]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux30~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~17 .lut_mask = 16'hF0CA;
defparam \Mux30~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N0
cycloneive_lcell_comb \Mux30~18 (
// Equation(s):
// \Mux30~18_combout  = (dcifimemload_22 & ((\Mux30~17_combout  & (\my_reg[15][1]~q )) # (!\Mux30~17_combout  & ((\my_reg[14][1]~q ))))) # (!dcifimemload_22 & (((\Mux30~17_combout ))))

	.dataa(\my_reg[15][1]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[14][1]~q ),
	.datad(\Mux30~17_combout ),
	.cin(gnd),
	.combout(\Mux30~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~18 .lut_mask = 16'hBBC0;
defparam \Mux30~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N23
dffeas \my_reg[31][31] (
	.clk(CLK),
	.d(wdat2),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][31] .is_wysiwyg = "true";
defparam \my_reg[31][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y36_N25
dffeas \my_reg[27][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][31] .is_wysiwyg = "true";
defparam \my_reg[27][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N8
cycloneive_lcell_comb \my_reg[19][31]~feeder (
// Equation(s):
// \my_reg[19][31]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat2),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[19][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[19][31]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[19][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N14
cycloneive_lcell_comb \Decoder0~29 (
// Equation(s):
// \Decoder0~29_combout  = (\wsel~4_combout  & (\wsel~2_combout  & (!\wsel~3_combout  & \Decoder0~12_combout )))

	.dataa(wsel4),
	.datab(wsel2),
	.datac(wsel3),
	.datad(\Decoder0~12_combout ),
	.cin(gnd),
	.combout(\Decoder0~29_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~29 .lut_mask = 16'h0800;
defparam \Decoder0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N9
dffeas \my_reg[19][31] (
	.clk(CLK),
	.d(\my_reg[19][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][31] .is_wysiwyg = "true";
defparam \my_reg[19][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N18
cycloneive_lcell_comb \Mux0~7 (
// Equation(s):
// \Mux0~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[23][31]~q )) # (!dcifimemload_23 & ((\my_reg[19][31]~q )))))

	.dataa(\my_reg[23][31]~q ),
	.datab(\my_reg[19][31]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~7 .lut_mask = 16'hFA0C;
defparam \Mux0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N24
cycloneive_lcell_comb \Mux0~8 (
// Equation(s):
// \Mux0~8_combout  = (dcifimemload_24 & ((\Mux0~7_combout  & (\my_reg[31][31]~q )) # (!\Mux0~7_combout  & ((\my_reg[27][31]~q ))))) # (!dcifimemload_24 & (((\Mux0~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[31][31]~q ),
	.datac(\my_reg[27][31]~q ),
	.datad(\Mux0~7_combout ),
	.cin(gnd),
	.combout(\Mux0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~8 .lut_mask = 16'hDDA0;
defparam \Mux0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N12
cycloneive_lcell_comb \my_reg[25][31]~feeder (
// Equation(s):
// \my_reg[25][31]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat2),
	.cin(gnd),
	.combout(\my_reg[25][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][31]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[25][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N13
dffeas \my_reg[25][31] (
	.clk(CLK),
	.d(\my_reg[25][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][31] .is_wysiwyg = "true";
defparam \my_reg[25][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N5
dffeas \my_reg[29][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][31] .is_wysiwyg = "true";
defparam \my_reg[29][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N30
cycloneive_lcell_comb \my_reg[21][31]~feeder (
// Equation(s):
// \my_reg[21][31]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat2),
	.cin(gnd),
	.combout(\my_reg[21][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][31]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[21][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N31
dffeas \my_reg[21][31] (
	.clk(CLK),
	.d(\my_reg[21][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][31] .is_wysiwyg = "true";
defparam \my_reg[21][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N0
cycloneive_lcell_comb \my_reg[17][31]~feeder (
// Equation(s):
// \my_reg[17][31]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat2),
	.cin(gnd),
	.combout(\my_reg[17][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[17][31]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[17][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N2
cycloneive_lcell_comb \Decoder0~14 (
// Equation(s):
// \Decoder0~14_combout  = (\wsel~0_combout  & (!\wsel~1_combout  & (\Decoder0~10_combout  & cuifRegWEN1)))

	.dataa(wsel),
	.datab(wsel1),
	.datac(\Decoder0~10_combout ),
	.datad(cuifRegWEN),
	.cin(gnd),
	.combout(\Decoder0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~14 .lut_mask = 16'h2000;
defparam \Decoder0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N1
dffeas \my_reg[17][31] (
	.clk(CLK),
	.d(\my_reg[17][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][31] .is_wysiwyg = "true";
defparam \my_reg[17][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N14
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// \Mux0~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[21][31]~q )) # (!dcifimemload_23 & ((\my_reg[17][31]~q )))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[21][31]~q ),
	.datac(\my_reg[17][31]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'hEE50;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N4
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// \Mux0~1_combout  = (dcifimemload_24 & ((\Mux0~0_combout  & ((\my_reg[29][31]~q ))) # (!\Mux0~0_combout  & (\my_reg[25][31]~q )))) # (!dcifimemload_24 & (((\Mux0~0_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[25][31]~q ),
	.datac(\my_reg[29][31]~q ),
	.datad(\Mux0~0_combout ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hF588;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N2
cycloneive_lcell_comb \Decoder0~25 (
// Equation(s):
// \Decoder0~25_combout  = (\wsel~3_combout  & (!\wsel~4_combout  & \Decoder0~19_combout ))

	.dataa(wsel3),
	.datab(gnd),
	.datac(wsel4),
	.datad(\Decoder0~19_combout ),
	.cin(gnd),
	.combout(\Decoder0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~25 .lut_mask = 16'h0A00;
defparam \Decoder0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N19
dffeas \my_reg[28][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][31] .is_wysiwyg = "true";
defparam \my_reg[28][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N1
dffeas \my_reg[20][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][31] .is_wysiwyg = "true";
defparam \my_reg[20][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N18
cycloneive_lcell_comb \Mux0~5 (
// Equation(s):
// \Mux0~5_combout  = (\Mux0~4_combout  & (((\my_reg[28][31]~q )) # (!dcifimemload_23))) # (!\Mux0~4_combout  & (dcifimemload_23 & ((\my_reg[20][31]~q ))))

	.dataa(\Mux0~4_combout ),
	.datab(dcifimemload_23),
	.datac(\my_reg[28][31]~q ),
	.datad(\my_reg[20][31]~q ),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~5 .lut_mask = 16'hE6A2;
defparam \Mux0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y42_N27
dffeas \my_reg[30][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][31] .is_wysiwyg = "true";
defparam \my_reg[30][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y42_N17
dffeas \my_reg[18][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][31] .is_wysiwyg = "true";
defparam \my_reg[18][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N16
cycloneive_lcell_comb \Mux0~2 (
// Equation(s):
// \Mux0~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[26][31]~q )) # (!dcifimemload_24 & ((\my_reg[18][31]~q )))))

	.dataa(\my_reg[26][31]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[18][31]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~2 .lut_mask = 16'hEE30;
defparam \Mux0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N26
cycloneive_lcell_comb \Mux0~3 (
// Equation(s):
// \Mux0~3_combout  = (dcifimemload_23 & ((\Mux0~2_combout  & ((\my_reg[30][31]~q ))) # (!\Mux0~2_combout  & (\my_reg[22][31]~q )))) # (!dcifimemload_23 & (((\Mux0~2_combout ))))

	.dataa(\my_reg[22][31]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[30][31]~q ),
	.datad(\Mux0~2_combout ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~3 .lut_mask = 16'hF388;
defparam \Mux0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N16
cycloneive_lcell_comb \Mux0~6 (
// Equation(s):
// \Mux0~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux0~3_combout ))) # (!dcifimemload_22 & (\Mux0~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux0~5_combout ),
	.datad(\Mux0~3_combout ),
	.cin(gnd),
	.combout(\Mux0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~6 .lut_mask = 16'hDC98;
defparam \Mux0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N26
cycloneive_lcell_comb \Mux0~9 (
// Equation(s):
// \Mux0~9_combout  = (dcifimemload_21 & ((\Mux0~6_combout  & (\Mux0~8_combout )) # (!\Mux0~6_combout  & ((\Mux0~1_combout ))))) # (!dcifimemload_21 & (((\Mux0~6_combout ))))

	.dataa(\Mux0~8_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux0~1_combout ),
	.datad(\Mux0~6_combout ),
	.cin(gnd),
	.combout(\Mux0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~9 .lut_mask = 16'hBBC0;
defparam \Mux0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y42_N11
dffeas \my_reg[9][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][31] .is_wysiwyg = "true";
defparam \my_reg[9][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N19
dffeas \my_reg[11][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][31] .is_wysiwyg = "true";
defparam \my_reg[11][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N25
dffeas \my_reg[8][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][31] .is_wysiwyg = "true";
defparam \my_reg[8][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N24
cycloneive_lcell_comb \Mux0~10 (
// Equation(s):
// \Mux0~10_combout  = (dcifimemload_22 & ((\my_reg[10][31]~q ) # ((dcifimemload_21)))) # (!dcifimemload_22 & (((\my_reg[8][31]~q  & !dcifimemload_21))))

	.dataa(\my_reg[10][31]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[8][31]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~10 .lut_mask = 16'hCCB8;
defparam \Mux0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N18
cycloneive_lcell_comb \Mux0~11 (
// Equation(s):
// \Mux0~11_combout  = (dcifimemload_21 & ((\Mux0~10_combout  & ((\my_reg[11][31]~q ))) # (!\Mux0~10_combout  & (\my_reg[9][31]~q )))) # (!dcifimemload_21 & (((\Mux0~10_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][31]~q ),
	.datac(\my_reg[11][31]~q ),
	.datad(\Mux0~10_combout ),
	.cin(gnd),
	.combout(\Mux0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~11 .lut_mask = 16'hF588;
defparam \Mux0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N23
dffeas \my_reg[15][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][31] .is_wysiwyg = "true";
defparam \my_reg[15][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N11
dffeas \my_reg[13][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][31] .is_wysiwyg = "true";
defparam \my_reg[13][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N25
dffeas \my_reg[12][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][31] .is_wysiwyg = "true";
defparam \my_reg[12][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N24
cycloneive_lcell_comb \Mux0~17 (
// Equation(s):
// \Mux0~17_combout  = (dcifimemload_21 & ((\my_reg[13][31]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][31]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[13][31]~q ),
	.datac(\my_reg[12][31]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~17 .lut_mask = 16'hAAD8;
defparam \Mux0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N22
cycloneive_lcell_comb \Mux0~18 (
// Equation(s):
// \Mux0~18_combout  = (dcifimemload_22 & ((\Mux0~17_combout  & ((\my_reg[15][31]~q ))) # (!\Mux0~17_combout  & (\my_reg[14][31]~q )))) # (!dcifimemload_22 & (((\Mux0~17_combout ))))

	.dataa(\my_reg[14][31]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[15][31]~q ),
	.datad(\Mux0~17_combout ),
	.cin(gnd),
	.combout(\Mux0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~18 .lut_mask = 16'hF388;
defparam \Mux0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y43_N15
dffeas \my_reg[2][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][31] .is_wysiwyg = "true";
defparam \my_reg[2][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y42_N13
dffeas \my_reg[3][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][31] .is_wysiwyg = "true";
defparam \my_reg[3][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y42_N15
dffeas \my_reg[1][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][31] .is_wysiwyg = "true";
defparam \my_reg[1][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N14
cycloneive_lcell_comb \Mux0~14 (
// Equation(s):
// \Mux0~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\my_reg[3][31]~q )) # (!dcifimemload_22 & ((\my_reg[1][31]~q )))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[3][31]~q ),
	.datac(\my_reg[1][31]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~14 .lut_mask = 16'h88A0;
defparam \Mux0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N14
cycloneive_lcell_comb \Mux0~15 (
// Equation(s):
// \Mux0~15_combout  = (\Mux0~14_combout ) # ((!dcifimemload_21 & (dcifimemload_22 & \my_reg[2][31]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\my_reg[2][31]~q ),
	.datad(\Mux0~14_combout ),
	.cin(gnd),
	.combout(\Mux0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~15 .lut_mask = 16'hFF40;
defparam \Mux0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y43_N21
dffeas \my_reg[7][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][31] .is_wysiwyg = "true";
defparam \my_reg[7][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N20
cycloneive_lcell_comb \my_reg[4][31]~feeder (
// Equation(s):
// \my_reg[4][31]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat2),
	.cin(gnd),
	.combout(\my_reg[4][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[4][31]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[4][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y43_N21
dffeas \my_reg[4][31] (
	.clk(CLK),
	.d(\my_reg[4][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][31] .is_wysiwyg = "true";
defparam \my_reg[4][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N18
cycloneive_lcell_comb \Mux0~12 (
// Equation(s):
// \Mux0~12_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\my_reg[5][31]~q )) # (!dcifimemload_21 & ((\my_reg[4][31]~q )))))

	.dataa(\my_reg[5][31]~q ),
	.datab(\my_reg[4][31]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~12 .lut_mask = 16'hFA0C;
defparam \Mux0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N20
cycloneive_lcell_comb \Mux0~13 (
// Equation(s):
// \Mux0~13_combout  = (dcifimemload_22 & ((\Mux0~12_combout  & ((\my_reg[7][31]~q ))) # (!\Mux0~12_combout  & (\my_reg[6][31]~q )))) # (!dcifimemload_22 & (((\Mux0~12_combout ))))

	.dataa(\my_reg[6][31]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[7][31]~q ),
	.datad(\Mux0~12_combout ),
	.cin(gnd),
	.combout(\Mux0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~13 .lut_mask = 16'hF388;
defparam \Mux0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N28
cycloneive_lcell_comb \Mux0~16 (
// Equation(s):
// \Mux0~16_combout  = (dcifimemload_23 & ((dcifimemload_24) # ((\Mux0~13_combout )))) # (!dcifimemload_23 & (!dcifimemload_24 & (\Mux0~15_combout )))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux0~15_combout ),
	.datad(\Mux0~13_combout ),
	.cin(gnd),
	.combout(\Mux0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~16 .lut_mask = 16'hBA98;
defparam \Mux0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N18
cycloneive_lcell_comb \Mux0~19 (
// Equation(s):
// \Mux0~19_combout  = (dcifimemload_24 & ((\Mux0~16_combout  & ((\Mux0~18_combout ))) # (!\Mux0~16_combout  & (\Mux0~11_combout )))) # (!dcifimemload_24 & (((\Mux0~16_combout ))))

	.dataa(dcifimemload_24),
	.datab(\Mux0~11_combout ),
	.datac(\Mux0~18_combout ),
	.datad(\Mux0~16_combout ),
	.cin(gnd),
	.combout(\Mux0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~19 .lut_mask = 16'hF588;
defparam \Mux0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N24
cycloneive_lcell_comb \my_reg[6][31]~feeder (
// Equation(s):
// \my_reg[6][31]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat2),
	.cin(gnd),
	.combout(\my_reg[6][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[6][31]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[6][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N25
dffeas \my_reg[6][31] (
	.clk(CLK),
	.d(\my_reg[6][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][31] .is_wysiwyg = "true";
defparam \my_reg[6][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N26
cycloneive_lcell_comb \Mux32~0 (
// Equation(s):
// \Mux32~0_combout  = (dcifimemload_16 & ((\my_reg[5][31]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\my_reg[4][31]~q  & !dcifimemload_17))))

	.dataa(\my_reg[5][31]~q ),
	.datab(\my_reg[4][31]~q ),
	.datac(dcifimemload_16),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux32~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~0 .lut_mask = 16'hF0AC;
defparam \Mux32~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N20
cycloneive_lcell_comb \Mux32~1 (
// Equation(s):
// \Mux32~1_combout  = (\Mux32~0_combout  & ((\my_reg[7][31]~q ) # ((!dcifimemload_17)))) # (!\Mux32~0_combout  & (((\my_reg[6][31]~q  & dcifimemload_17))))

	.dataa(\my_reg[7][31]~q ),
	.datab(\my_reg[6][31]~q ),
	.datac(\Mux32~0_combout ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux32~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~1 .lut_mask = 16'hACF0;
defparam \Mux32~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N16
cycloneive_lcell_comb \my_reg[14][31]~feeder (
// Equation(s):
// \my_reg[14][31]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat2),
	.cin(gnd),
	.combout(\my_reg[14][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[14][31]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[14][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N17
dffeas \my_reg[14][31] (
	.clk(CLK),
	.d(\my_reg[14][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][31] .is_wysiwyg = "true";
defparam \my_reg[14][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N10
cycloneive_lcell_comb \Mux32~7 (
// Equation(s):
// \Mux32~7_combout  = (dcifimemload_16 & (((\my_reg[13][31]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[12][31]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[12][31]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[13][31]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux32~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~7 .lut_mask = 16'hCCE2;
defparam \Mux32~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N24
cycloneive_lcell_comb \Mux32~8 (
// Equation(s):
// \Mux32~8_combout  = (dcifimemload_17 & ((\Mux32~7_combout  & ((\my_reg[15][31]~q ))) # (!\Mux32~7_combout  & (\my_reg[14][31]~q )))) # (!dcifimemload_17 & (((\Mux32~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[14][31]~q ),
	.datac(\my_reg[15][31]~q ),
	.datad(\Mux32~7_combout ),
	.cin(gnd),
	.combout(\Mux32~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~8 .lut_mask = 16'hF588;
defparam \Mux32~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N10
cycloneive_lcell_comb \Mux32~3 (
// Equation(s):
// \Mux32~3_combout  = (\Mux32~2_combout  & ((\my_reg[11][31]~q ) # ((!dcifimemload_16)))) # (!\Mux32~2_combout  & (((\my_reg[9][31]~q  & dcifimemload_16))))

	.dataa(\Mux32~2_combout ),
	.datab(\my_reg[11][31]~q ),
	.datac(\my_reg[9][31]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux32~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~3 .lut_mask = 16'hD8AA;
defparam \Mux32~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N12
cycloneive_lcell_comb \Mux32~4 (
// Equation(s):
// \Mux32~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][31]~q ))) # (!dcifimemload_17 & (\my_reg[1][31]~q ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[1][31]~q ),
	.datac(\my_reg[3][31]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux32~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~4 .lut_mask = 16'hA088;
defparam \Mux32~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N18
cycloneive_lcell_comb \Mux32~5 (
// Equation(s):
// \Mux32~5_combout  = (\Mux32~4_combout ) # ((!dcifimemload_16 & (\my_reg[2][31]~q  & dcifimemload_17)))

	.dataa(dcifimemload_16),
	.datab(\my_reg[2][31]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux32~4_combout ),
	.cin(gnd),
	.combout(\Mux32~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~5 .lut_mask = 16'hFF40;
defparam \Mux32~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N28
cycloneive_lcell_comb \Mux32~6 (
// Equation(s):
// \Mux32~6_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\Mux32~3_combout )))) # (!dcifimemload_19 & (!dcifimemload_18 & ((\Mux32~5_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux32~3_combout ),
	.datad(\Mux32~5_combout ),
	.cin(gnd),
	.combout(\Mux32~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~6 .lut_mask = 16'hB9A8;
defparam \Mux32~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N8
cycloneive_lcell_comb \my_reg[23][31]~feeder (
// Equation(s):
// \my_reg[23][31]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat2),
	.cin(gnd),
	.combout(\my_reg[23][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[23][31]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[23][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N9
dffeas \my_reg[23][31] (
	.clk(CLK),
	.d(\my_reg[23][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][31] .is_wysiwyg = "true";
defparam \my_reg[23][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N2
cycloneive_lcell_comb \Mux32~17 (
// Equation(s):
// \Mux32~17_combout  = (dcifimemload_19 & (((\my_reg[27][31]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[19][31]~q  & ((!dcifimemload_18))))

	.dataa(\my_reg[19][31]~q ),
	.datab(\my_reg[27][31]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux32~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~17 .lut_mask = 16'hF0CA;
defparam \Mux32~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N20
cycloneive_lcell_comb \Mux32~18 (
// Equation(s):
// \Mux32~18_combout  = (dcifimemload_18 & ((\Mux32~17_combout  & (\my_reg[31][31]~q )) # (!\Mux32~17_combout  & ((\my_reg[23][31]~q ))))) # (!dcifimemload_18 & (((\Mux32~17_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[31][31]~q ),
	.datac(\my_reg[23][31]~q ),
	.datad(\Mux32~17_combout ),
	.cin(gnd),
	.combout(\Mux32~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~18 .lut_mask = 16'hDDA0;
defparam \Mux32~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N28
cycloneive_lcell_comb \Mux32~10 (
// Equation(s):
// \Mux32~10_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[25][31]~q ))) # (!dcifimemload_19 & (\my_reg[17][31]~q ))))

	.dataa(\my_reg[17][31]~q ),
	.datab(\my_reg[25][31]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux32~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~10 .lut_mask = 16'hFC0A;
defparam \Mux32~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N2
cycloneive_lcell_comb \Mux32~11 (
// Equation(s):
// \Mux32~11_combout  = (dcifimemload_18 & ((\Mux32~10_combout  & ((\my_reg[29][31]~q ))) # (!\Mux32~10_combout  & (\my_reg[21][31]~q )))) # (!dcifimemload_18 & (((\Mux32~10_combout ))))

	.dataa(\my_reg[21][31]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[29][31]~q ),
	.datad(\Mux32~10_combout ),
	.cin(gnd),
	.combout(\Mux32~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~11 .lut_mask = 16'hF388;
defparam \Mux32~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N31
dffeas \my_reg[24][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][31] .is_wysiwyg = "true";
defparam \my_reg[24][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N13
dffeas \my_reg[16][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][31] .is_wysiwyg = "true";
defparam \my_reg[16][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N0
cycloneive_lcell_comb \Mux32~14 (
// Equation(s):
// \Mux32~14_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[20][31]~q ))) # (!dcifimemload_18 & (\my_reg[16][31]~q ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[16][31]~q ),
	.datac(\my_reg[20][31]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux32~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~14 .lut_mask = 16'hFA44;
defparam \Mux32~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N30
cycloneive_lcell_comb \Mux32~15 (
// Equation(s):
// \Mux32~15_combout  = (dcifimemload_19 & ((\Mux32~14_combout  & (\my_reg[28][31]~q )) # (!\Mux32~14_combout  & ((\my_reg[24][31]~q ))))) # (!dcifimemload_19 & (((\Mux32~14_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[28][31]~q ),
	.datac(\my_reg[24][31]~q ),
	.datad(\Mux32~14_combout ),
	.cin(gnd),
	.combout(\Mux32~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~15 .lut_mask = 16'hDDA0;
defparam \Mux32~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N19
dffeas \my_reg[26][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][31] .is_wysiwyg = "true";
defparam \my_reg[26][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N0
cycloneive_lcell_comb \Decoder0~18 (
// Equation(s):
// \Decoder0~18_combout  = (\wsel~3_combout  & (\wsel~4_combout  & \Decoder0~17_combout ))

	.dataa(wsel3),
	.datab(gnd),
	.datac(wsel4),
	.datad(\Decoder0~17_combout ),
	.cin(gnd),
	.combout(\Decoder0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~18 .lut_mask = 16'hA000;
defparam \Decoder0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N17
dffeas \my_reg[22][31] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][31] .is_wysiwyg = "true";
defparam \my_reg[22][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N16
cycloneive_lcell_comb \Mux32~12 (
// Equation(s):
// \Mux32~12_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[22][31]~q ))) # (!dcifimemload_18 & (\my_reg[18][31]~q ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[18][31]~q ),
	.datac(\my_reg[22][31]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux32~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~12 .lut_mask = 16'hFA44;
defparam \Mux32~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N18
cycloneive_lcell_comb \Mux32~13 (
// Equation(s):
// \Mux32~13_combout  = (dcifimemload_19 & ((\Mux32~12_combout  & (\my_reg[30][31]~q )) # (!\Mux32~12_combout  & ((\my_reg[26][31]~q ))))) # (!dcifimemload_19 & (((\Mux32~12_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[30][31]~q ),
	.datac(\my_reg[26][31]~q ),
	.datad(\Mux32~12_combout ),
	.cin(gnd),
	.combout(\Mux32~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~13 .lut_mask = 16'hDDA0;
defparam \Mux32~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N2
cycloneive_lcell_comb \Mux32~16 (
// Equation(s):
// \Mux32~16_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux32~13_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & (\Mux32~15_combout )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux32~15_combout ),
	.datad(\Mux32~13_combout ),
	.cin(gnd),
	.combout(\Mux32~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~16 .lut_mask = 16'hBA98;
defparam \Mux32~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N7
dffeas \my_reg[31][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][30] .is_wysiwyg = "true";
defparam \my_reg[31][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N29
dffeas \my_reg[19][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][30] .is_wysiwyg = "true";
defparam \my_reg[19][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N28
cycloneive_lcell_comb \Mux1~7 (
// Equation(s):
// \Mux1~7_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[27][30]~q )) # (!dcifimemload_24 & ((\my_reg[19][30]~q )))))

	.dataa(\my_reg[27][30]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[19][30]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux1~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~7 .lut_mask = 16'hEE30;
defparam \Mux1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N6
cycloneive_lcell_comb \Mux1~8 (
// Equation(s):
// \Mux1~8_combout  = (dcifimemload_23 & ((\Mux1~7_combout  & ((\my_reg[31][30]~q ))) # (!\Mux1~7_combout  & (\my_reg[23][30]~q )))) # (!dcifimemload_23 & (((\Mux1~7_combout ))))

	.dataa(\my_reg[23][30]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[31][30]~q ),
	.datad(\Mux1~7_combout ),
	.cin(gnd),
	.combout(\Mux1~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~8 .lut_mask = 16'hF388;
defparam \Mux1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N15
dffeas \my_reg[22][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][30] .is_wysiwyg = "true";
defparam \my_reg[22][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N9
dffeas \my_reg[18][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][30] .is_wysiwyg = "true";
defparam \my_reg[18][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N8
cycloneive_lcell_comb \Mux1~2 (
// Equation(s):
// \Mux1~2_combout  = (dcifimemload_23 & ((\my_reg[22][30]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[18][30]~q  & !dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[22][30]~q ),
	.datac(\my_reg[18][30]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~2 .lut_mask = 16'hAAD8;
defparam \Mux1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N3
dffeas \my_reg[30][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][30] .is_wysiwyg = "true";
defparam \my_reg[30][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N2
cycloneive_lcell_comb \Mux1~3 (
// Equation(s):
// \Mux1~3_combout  = (\Mux1~2_combout  & (((\my_reg[30][30]~q ) # (!dcifimemload_24)))) # (!\Mux1~2_combout  & (\my_reg[26][30]~q  & ((dcifimemload_24))))

	.dataa(\my_reg[26][30]~q ),
	.datab(\Mux1~2_combout ),
	.datac(\my_reg[30][30]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~3 .lut_mask = 16'hE2CC;
defparam \Mux1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y40_N1
dffeas \my_reg[24][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][30] .is_wysiwyg = "true";
defparam \my_reg[24][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N15
dffeas \my_reg[28][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][30] .is_wysiwyg = "true";
defparam \my_reg[28][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N31
dffeas \my_reg[20][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][30] .is_wysiwyg = "true";
defparam \my_reg[20][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N21
dffeas \my_reg[16][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][30] .is_wysiwyg = "true";
defparam \my_reg[16][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N20
cycloneive_lcell_comb \Mux1~4 (
// Equation(s):
// \Mux1~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[20][30]~q )) # (!dcifimemload_23 & ((\my_reg[16][30]~q )))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[20][30]~q ),
	.datac(\my_reg[16][30]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~4 .lut_mask = 16'hEE50;
defparam \Mux1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N14
cycloneive_lcell_comb \Mux1~5 (
// Equation(s):
// \Mux1~5_combout  = (dcifimemload_24 & ((\Mux1~4_combout  & ((\my_reg[28][30]~q ))) # (!\Mux1~4_combout  & (\my_reg[24][30]~q )))) # (!dcifimemload_24 & (((\Mux1~4_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[24][30]~q ),
	.datac(\my_reg[28][30]~q ),
	.datad(\Mux1~4_combout ),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~5 .lut_mask = 16'hF588;
defparam \Mux1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N4
cycloneive_lcell_comb \Mux1~6 (
// Equation(s):
// \Mux1~6_combout  = (dcifimemload_22 & ((\Mux1~3_combout ) # ((dcifimemload_21)))) # (!dcifimemload_22 & (((\Mux1~5_combout  & !dcifimemload_21))))

	.dataa(dcifimemload_22),
	.datab(\Mux1~3_combout ),
	.datac(\Mux1~5_combout ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux1~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~6 .lut_mask = 16'hAAD8;
defparam \Mux1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N0
cycloneive_lcell_comb \my_reg[21][30]~feeder (
// Equation(s):
// \my_reg[21][30]~feeder_combout  = \wdat~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat3),
	.cin(gnd),
	.combout(\my_reg[21][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][30]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[21][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N1
dffeas \my_reg[21][30] (
	.clk(CLK),
	.d(\my_reg[21][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][30] .is_wysiwyg = "true";
defparam \my_reg[21][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N15
dffeas \my_reg[29][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][30] .is_wysiwyg = "true";
defparam \my_reg[29][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N30
cycloneive_lcell_comb \my_reg[25][30]~feeder (
// Equation(s):
// \my_reg[25][30]~feeder_combout  = \wdat~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat3),
	.cin(gnd),
	.combout(\my_reg[25][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][30]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[25][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N31
dffeas \my_reg[25][30] (
	.clk(CLK),
	.d(\my_reg[25][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][30] .is_wysiwyg = "true";
defparam \my_reg[25][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N23
dffeas \my_reg[17][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][30] .is_wysiwyg = "true";
defparam \my_reg[17][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N22
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[25][30]~q )) # (!dcifimemload_24 & ((\my_reg[17][30]~q )))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[25][30]~q ),
	.datac(\my_reg[17][30]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'hEE50;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N14
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// \Mux1~1_combout  = (dcifimemload_23 & ((\Mux1~0_combout  & ((\my_reg[29][30]~q ))) # (!\Mux1~0_combout  & (\my_reg[21][30]~q )))) # (!dcifimemload_23 & (((\Mux1~0_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[21][30]~q ),
	.datac(\my_reg[29][30]~q ),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hF588;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N14
cycloneive_lcell_comb \Mux1~9 (
// Equation(s):
// \Mux1~9_combout  = (dcifimemload_21 & ((\Mux1~6_combout  & (\Mux1~8_combout )) # (!\Mux1~6_combout  & ((\Mux1~1_combout ))))) # (!dcifimemload_21 & (((\Mux1~6_combout ))))

	.dataa(\Mux1~8_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux1~6_combout ),
	.datad(\Mux1~1_combout ),
	.cin(gnd),
	.combout(\Mux1~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~9 .lut_mask = 16'hBCB0;
defparam \Mux1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N3
dffeas \my_reg[9][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][30] .is_wysiwyg = "true";
defparam \my_reg[9][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N31
dffeas \my_reg[11][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][30] .is_wysiwyg = "true";
defparam \my_reg[11][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N13
dffeas \my_reg[8][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][30] .is_wysiwyg = "true";
defparam \my_reg[8][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N12
cycloneive_lcell_comb \Mux1~12 (
// Equation(s):
// \Mux1~12_combout  = (dcifimemload_22 & ((\my_reg[10][30]~q ) # ((dcifimemload_21)))) # (!dcifimemload_22 & (((\my_reg[8][30]~q  & !dcifimemload_21))))

	.dataa(\my_reg[10][30]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[8][30]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux1~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~12 .lut_mask = 16'hCCB8;
defparam \Mux1~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N30
cycloneive_lcell_comb \Mux1~13 (
// Equation(s):
// \Mux1~13_combout  = (dcifimemload_21 & ((\Mux1~12_combout  & ((\my_reg[11][30]~q ))) # (!\Mux1~12_combout  & (\my_reg[9][30]~q )))) # (!dcifimemload_21 & (((\Mux1~12_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][30]~q ),
	.datac(\my_reg[11][30]~q ),
	.datad(\Mux1~12_combout ),
	.cin(gnd),
	.combout(\Mux1~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~13 .lut_mask = 16'hF588;
defparam \Mux1~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N16
cycloneive_lcell_comb \my_reg[2][30]~feeder (
// Equation(s):
// \my_reg[2][30]~feeder_combout  = \wdat~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat3),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[2][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[2][30]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[2][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N17
dffeas \my_reg[2][30] (
	.clk(CLK),
	.d(\my_reg[2][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][30] .is_wysiwyg = "true";
defparam \my_reg[2][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y42_N7
dffeas \my_reg[1][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][30] .is_wysiwyg = "true";
defparam \my_reg[1][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y42_N25
dffeas \my_reg[3][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][30] .is_wysiwyg = "true";
defparam \my_reg[3][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N6
cycloneive_lcell_comb \Mux1~14 (
// Equation(s):
// \Mux1~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][30]~q ))) # (!dcifimemload_22 & (\my_reg[1][30]~q ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\my_reg[1][30]~q ),
	.datad(\my_reg[3][30]~q ),
	.cin(gnd),
	.combout(\Mux1~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~14 .lut_mask = 16'hA820;
defparam \Mux1~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N20
cycloneive_lcell_comb \Mux1~15 (
// Equation(s):
// \Mux1~15_combout  = (\Mux1~14_combout ) # ((dcifimemload_22 & (\my_reg[2][30]~q  & !dcifimemload_21)))

	.dataa(dcifimemload_22),
	.datab(\my_reg[2][30]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux1~14_combout ),
	.cin(gnd),
	.combout(\Mux1~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~15 .lut_mask = 16'hFF08;
defparam \Mux1~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N0
cycloneive_lcell_comb \Mux1~16 (
// Equation(s):
// \Mux1~16_combout  = (dcifimemload_24 & ((dcifimemload_23) # ((\Mux1~13_combout )))) # (!dcifimemload_24 & (!dcifimemload_23 & ((\Mux1~15_combout ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux1~13_combout ),
	.datad(\Mux1~15_combout ),
	.cin(gnd),
	.combout(\Mux1~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~16 .lut_mask = 16'hB9A8;
defparam \Mux1~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N3
dffeas \my_reg[15][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][30] .is_wysiwyg = "true";
defparam \my_reg[15][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N0
cycloneive_lcell_comb \my_reg[13][30]~feeder (
// Equation(s):
// \my_reg[13][30]~feeder_combout  = \wdat~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat3),
	.cin(gnd),
	.combout(\my_reg[13][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[13][30]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[13][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N1
dffeas \my_reg[13][30] (
	.clk(CLK),
	.d(\my_reg[13][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][30] .is_wysiwyg = "true";
defparam \my_reg[13][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N23
dffeas \my_reg[12][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][30] .is_wysiwyg = "true";
defparam \my_reg[12][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N22
cycloneive_lcell_comb \Mux1~17 (
// Equation(s):
// \Mux1~17_combout  = (dcifimemload_21 & ((\my_reg[13][30]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][30]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[13][30]~q ),
	.datac(\my_reg[12][30]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux1~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~17 .lut_mask = 16'hAAD8;
defparam \Mux1~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N2
cycloneive_lcell_comb \Mux1~18 (
// Equation(s):
// \Mux1~18_combout  = (dcifimemload_22 & ((\Mux1~17_combout  & ((\my_reg[15][30]~q ))) # (!\Mux1~17_combout  & (\my_reg[14][30]~q )))) # (!dcifimemload_22 & (((\Mux1~17_combout ))))

	.dataa(\my_reg[14][30]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[15][30]~q ),
	.datad(\Mux1~17_combout ),
	.cin(gnd),
	.combout(\Mux1~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~18 .lut_mask = 16'hF388;
defparam \Mux1~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N28
cycloneive_lcell_comb \my_reg[6][30]~feeder (
// Equation(s):
// \my_reg[6][30]~feeder_combout  = \wdat~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat3),
	.cin(gnd),
	.combout(\my_reg[6][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[6][30]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[6][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N29
dffeas \my_reg[6][30] (
	.clk(CLK),
	.d(\my_reg[6][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][30] .is_wysiwyg = "true";
defparam \my_reg[6][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N3
dffeas \my_reg[7][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][30] .is_wysiwyg = "true";
defparam \my_reg[7][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N24
cycloneive_lcell_comb \my_reg[5][30]~feeder (
// Equation(s):
// \my_reg[5][30]~feeder_combout  = \wdat~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat3),
	.cin(gnd),
	.combout(\my_reg[5][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[5][30]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[5][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y38_N25
dffeas \my_reg[5][30] (
	.clk(CLK),
	.d(\my_reg[5][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][30] .is_wysiwyg = "true";
defparam \my_reg[5][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N30
cycloneive_lcell_comb \Mux1~10 (
// Equation(s):
// \Mux1~10_combout  = (dcifimemload_21 & (((\my_reg[5][30]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\my_reg[4][30]~q  & ((!dcifimemload_22))))

	.dataa(\my_reg[4][30]~q ),
	.datab(\my_reg[5][30]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~10 .lut_mask = 16'hF0CA;
defparam \Mux1~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N22
cycloneive_lcell_comb \Mux1~11 (
// Equation(s):
// \Mux1~11_combout  = (dcifimemload_22 & ((\Mux1~10_combout  & ((\my_reg[7][30]~q ))) # (!\Mux1~10_combout  & (\my_reg[6][30]~q )))) # (!dcifimemload_22 & (((\Mux1~10_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[6][30]~q ),
	.datac(\my_reg[7][30]~q ),
	.datad(\Mux1~10_combout ),
	.cin(gnd),
	.combout(\Mux1~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~11 .lut_mask = 16'hF588;
defparam \Mux1~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N6
cycloneive_lcell_comb \Mux1~19 (
// Equation(s):
// \Mux1~19_combout  = (dcifimemload_23 & ((\Mux1~16_combout  & (\Mux1~18_combout )) # (!\Mux1~16_combout  & ((\Mux1~11_combout ))))) # (!dcifimemload_23 & (\Mux1~16_combout ))

	.dataa(dcifimemload_23),
	.datab(\Mux1~16_combout ),
	.datac(\Mux1~18_combout ),
	.datad(\Mux1~11_combout ),
	.cin(gnd),
	.combout(\Mux1~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~19 .lut_mask = 16'hE6C4;
defparam \Mux1~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N14
cycloneive_lcell_comb \Mux33~0 (
// Equation(s):
// \Mux33~0_combout  = (dcifimemload_17 & ((\my_reg[10][30]~q ) # ((dcifimemload_16)))) # (!dcifimemload_17 & (((\my_reg[8][30]~q  & !dcifimemload_16))))

	.dataa(\my_reg[10][30]~q ),
	.datab(dcifimemload_17),
	.datac(\my_reg[8][30]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux33~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~0 .lut_mask = 16'hCCB8;
defparam \Mux33~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N16
cycloneive_lcell_comb \Mux33~1 (
// Equation(s):
// \Mux33~1_combout  = (dcifimemload_16 & ((\Mux33~0_combout  & (\my_reg[11][30]~q )) # (!\Mux33~0_combout  & ((\my_reg[9][30]~q ))))) # (!dcifimemload_16 & (((\Mux33~0_combout ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[11][30]~q ),
	.datac(\my_reg[9][30]~q ),
	.datad(\Mux33~0_combout ),
	.cin(gnd),
	.combout(\Mux33~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~1 .lut_mask = 16'hDDA0;
defparam \Mux33~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N21
dffeas \my_reg[4][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][30] .is_wysiwyg = "true";
defparam \my_reg[4][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N20
cycloneive_lcell_comb \Mux33~2 (
// Equation(s):
// \Mux33~2_combout  = (dcifimemload_16 & ((\my_reg[5][30]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\my_reg[4][30]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[5][30]~q ),
	.datac(\my_reg[4][30]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux33~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~2 .lut_mask = 16'hAAD8;
defparam \Mux33~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N2
cycloneive_lcell_comb \Mux33~3 (
// Equation(s):
// \Mux33~3_combout  = (dcifimemload_17 & ((\Mux33~2_combout  & ((\my_reg[7][30]~q ))) # (!\Mux33~2_combout  & (\my_reg[6][30]~q )))) # (!dcifimemload_17 & (((\Mux33~2_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[6][30]~q ),
	.datac(\my_reg[7][30]~q ),
	.datad(\Mux33~2_combout ),
	.cin(gnd),
	.combout(\Mux33~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~3 .lut_mask = 16'hF588;
defparam \Mux33~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N24
cycloneive_lcell_comb \Mux33~4 (
// Equation(s):
// \Mux33~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][30]~q ))) # (!dcifimemload_17 & (\my_reg[1][30]~q ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[1][30]~q ),
	.datac(\my_reg[3][30]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux33~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~4 .lut_mask = 16'hA088;
defparam \Mux33~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N26
cycloneive_lcell_comb \Mux33~5 (
// Equation(s):
// \Mux33~5_combout  = (\Mux33~4_combout ) # ((!dcifimemload_16 & (\my_reg[2][30]~q  & dcifimemload_17)))

	.dataa(dcifimemload_16),
	.datab(\my_reg[2][30]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux33~4_combout ),
	.cin(gnd),
	.combout(\Mux33~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~5 .lut_mask = 16'hFF40;
defparam \Mux33~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N22
cycloneive_lcell_comb \Mux33~6 (
// Equation(s):
// \Mux33~6_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & (\Mux33~3_combout )) # (!dcifimemload_18 & ((\Mux33~5_combout )))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux33~3_combout ),
	.datad(\Mux33~5_combout ),
	.cin(gnd),
	.combout(\Mux33~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~6 .lut_mask = 16'hD9C8;
defparam \Mux33~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N9
dffeas \my_reg[14][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][30] .is_wysiwyg = "true";
defparam \my_reg[14][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N30
cycloneive_lcell_comb \Mux33~7 (
// Equation(s):
// \Mux33~7_combout  = (dcifimemload_16 & (((\my_reg[13][30]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[12][30]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[12][30]~q ),
	.datab(\my_reg[13][30]~q ),
	.datac(dcifimemload_16),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux33~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~7 .lut_mask = 16'hF0CA;
defparam \Mux33~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N8
cycloneive_lcell_comb \Mux33~8 (
// Equation(s):
// \Mux33~8_combout  = (dcifimemload_17 & ((\Mux33~7_combout  & (\my_reg[15][30]~q )) # (!\Mux33~7_combout  & ((\my_reg[14][30]~q ))))) # (!dcifimemload_17 & (((\Mux33~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[15][30]~q ),
	.datac(\my_reg[14][30]~q ),
	.datad(\Mux33~7_combout ),
	.cin(gnd),
	.combout(\Mux33~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~8 .lut_mask = 16'hDDA0;
defparam \Mux33~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N8
cycloneive_lcell_comb \Mux33~10 (
// Equation(s):
// \Mux33~10_combout  = (dcifimemload_18 & (((\my_reg[21][30]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[17][30]~q  & ((!dcifimemload_19))))

	.dataa(\my_reg[17][30]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[21][30]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux33~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~10 .lut_mask = 16'hCCE2;
defparam \Mux33~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N14
cycloneive_lcell_comb \Mux33~11 (
// Equation(s):
// \Mux33~11_combout  = (\Mux33~10_combout  & (((\my_reg[29][30]~q ) # (!dcifimemload_19)))) # (!\Mux33~10_combout  & (\my_reg[25][30]~q  & ((dcifimemload_19))))

	.dataa(\my_reg[25][30]~q ),
	.datab(\my_reg[29][30]~q ),
	.datac(\Mux33~10_combout ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux33~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~11 .lut_mask = 16'hCAF0;
defparam \Mux33~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N19
dffeas \my_reg[27][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][30] .is_wysiwyg = "true";
defparam \my_reg[27][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N15
dffeas \my_reg[23][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][30] .is_wysiwyg = "true";
defparam \my_reg[23][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N14
cycloneive_lcell_comb \Mux33~17 (
// Equation(s):
// \Mux33~17_combout  = (dcifimemload_18 & (((\my_reg[23][30]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[19][30]~q  & ((!dcifimemload_19))))

	.dataa(\my_reg[19][30]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[23][30]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux33~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~17 .lut_mask = 16'hCCE2;
defparam \Mux33~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N24
cycloneive_lcell_comb \Mux33~18 (
// Equation(s):
// \Mux33~18_combout  = (dcifimemload_19 & ((\Mux33~17_combout  & (\my_reg[31][30]~q )) # (!\Mux33~17_combout  & ((\my_reg[27][30]~q ))))) # (!dcifimemload_19 & (((\Mux33~17_combout ))))

	.dataa(\my_reg[31][30]~q ),
	.datab(\my_reg[27][30]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux33~17_combout ),
	.cin(gnd),
	.combout(\Mux33~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~18 .lut_mask = 16'hAFC0;
defparam \Mux33~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N0
cycloneive_lcell_comb \Mux33~14 (
// Equation(s):
// \Mux33~14_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & (\my_reg[24][30]~q )) # (!dcifimemload_19 & ((\my_reg[16][30]~q )))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\my_reg[24][30]~q ),
	.datad(\my_reg[16][30]~q ),
	.cin(gnd),
	.combout(\Mux33~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~14 .lut_mask = 16'hD9C8;
defparam \Mux33~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N30
cycloneive_lcell_comb \Mux33~15 (
// Equation(s):
// \Mux33~15_combout  = (dcifimemload_18 & ((\Mux33~14_combout  & (\my_reg[28][30]~q )) # (!\Mux33~14_combout  & ((\my_reg[20][30]~q ))))) # (!dcifimemload_18 & (((\Mux33~14_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[28][30]~q ),
	.datac(\my_reg[20][30]~q ),
	.datad(\Mux33~14_combout ),
	.cin(gnd),
	.combout(\Mux33~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~15 .lut_mask = 16'hDDA0;
defparam \Mux33~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N13
dffeas \my_reg[26][30] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][30] .is_wysiwyg = "true";
defparam \my_reg[26][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N12
cycloneive_lcell_comb \Mux33~12 (
// Equation(s):
// \Mux33~12_combout  = (dcifimemload_19 & (((\my_reg[26][30]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[18][30]~q  & ((!dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[18][30]~q ),
	.datac(\my_reg[26][30]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux33~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~12 .lut_mask = 16'hAAE4;
defparam \Mux33~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N14
cycloneive_lcell_comb \Mux33~13 (
// Equation(s):
// \Mux33~13_combout  = (dcifimemload_18 & ((\Mux33~12_combout  & (\my_reg[30][30]~q )) # (!\Mux33~12_combout  & ((\my_reg[22][30]~q ))))) # (!dcifimemload_18 & (((\Mux33~12_combout ))))

	.dataa(\my_reg[30][30]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[22][30]~q ),
	.datad(\Mux33~12_combout ),
	.cin(gnd),
	.combout(\Mux33~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~13 .lut_mask = 16'hBBC0;
defparam \Mux33~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N24
cycloneive_lcell_comb \Mux33~16 (
// Equation(s):
// \Mux33~16_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux33~13_combout ))) # (!dcifimemload_17 & (\Mux33~15_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux33~15_combout ),
	.datad(\Mux33~13_combout ),
	.cin(gnd),
	.combout(\Mux33~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~16 .lut_mask = 16'hDC98;
defparam \Mux33~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N25
dffeas \my_reg[6][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][29] .is_wysiwyg = "true";
defparam \my_reg[6][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N21
dffeas \my_reg[7][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][29] .is_wysiwyg = "true";
defparam \my_reg[7][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y42_N15
dffeas \my_reg[5][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][29] .is_wysiwyg = "true";
defparam \my_reg[5][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N11
dffeas \my_reg[4][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][29] .is_wysiwyg = "true";
defparam \my_reg[4][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N10
cycloneive_lcell_comb \Mux2~12 (
// Equation(s):
// \Mux2~12_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\my_reg[5][29]~q )) # (!dcifimemload_21 & ((\my_reg[4][29]~q )))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[5][29]~q ),
	.datac(\my_reg[4][29]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~12 .lut_mask = 16'hEE50;
defparam \Mux2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N20
cycloneive_lcell_comb \Mux2~13 (
// Equation(s):
// \Mux2~13_combout  = (dcifimemload_22 & ((\Mux2~12_combout  & ((\my_reg[7][29]~q ))) # (!\Mux2~12_combout  & (\my_reg[6][29]~q )))) # (!dcifimemload_22 & (((\Mux2~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[6][29]~q ),
	.datac(\my_reg[7][29]~q ),
	.datad(\Mux2~12_combout ),
	.cin(gnd),
	.combout(\Mux2~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~13 .lut_mask = 16'hF588;
defparam \Mux2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y43_N11
dffeas \my_reg[2][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][29] .is_wysiwyg = "true";
defparam \my_reg[2][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y42_N29
dffeas \my_reg[3][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][29] .is_wysiwyg = "true";
defparam \my_reg[3][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N0
cycloneive_lcell_comb \Mux2~14 (
// Equation(s):
// \Mux2~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][29]~q ))) # (!dcifimemload_22 & (\my_reg[1][29]~q ))))

	.dataa(\my_reg[1][29]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[3][29]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux2~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~14 .lut_mask = 16'hE200;
defparam \Mux2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N10
cycloneive_lcell_comb \Mux2~15 (
// Equation(s):
// \Mux2~15_combout  = (\Mux2~14_combout ) # ((!dcifimemload_21 & (dcifimemload_22 & \my_reg[2][29]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\my_reg[2][29]~q ),
	.datad(\Mux2~14_combout ),
	.cin(gnd),
	.combout(\Mux2~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~15 .lut_mask = 16'hFF40;
defparam \Mux2~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N10
cycloneive_lcell_comb \Mux2~16 (
// Equation(s):
// \Mux2~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & (\Mux2~13_combout )) # (!dcifimemload_23 & ((\Mux2~15_combout )))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux2~13_combout ),
	.datad(\Mux2~15_combout ),
	.cin(gnd),
	.combout(\Mux2~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~16 .lut_mask = 16'hD9C8;
defparam \Mux2~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y42_N25
dffeas \my_reg[10][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][29] .is_wysiwyg = "true";
defparam \my_reg[10][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N1
dffeas \my_reg[8][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][29] .is_wysiwyg = "true";
defparam \my_reg[8][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N0
cycloneive_lcell_comb \Mux2~10 (
// Equation(s):
// \Mux2~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][29]~q )) # (!dcifimemload_22 & ((\my_reg[8][29]~q )))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[10][29]~q ),
	.datac(\my_reg[8][29]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~10 .lut_mask = 16'hEE50;
defparam \Mux2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N27
dffeas \my_reg[11][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][29] .is_wysiwyg = "true";
defparam \my_reg[11][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N26
cycloneive_lcell_comb \Mux2~11 (
// Equation(s):
// \Mux2~11_combout  = (\Mux2~10_combout  & (((\my_reg[11][29]~q ) # (!dcifimemload_21)))) # (!\Mux2~10_combout  & (\my_reg[9][29]~q  & ((dcifimemload_21))))

	.dataa(\my_reg[9][29]~q ),
	.datab(\Mux2~10_combout ),
	.datac(\my_reg[11][29]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~11 .lut_mask = 16'hE2CC;
defparam \Mux2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N19
dffeas \my_reg[15][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][29] .is_wysiwyg = "true";
defparam \my_reg[15][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N23
dffeas \my_reg[13][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][29] .is_wysiwyg = "true";
defparam \my_reg[13][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N5
dffeas \my_reg[12][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][29] .is_wysiwyg = "true";
defparam \my_reg[12][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N4
cycloneive_lcell_comb \Mux2~17 (
// Equation(s):
// \Mux2~17_combout  = (dcifimemload_21 & ((\my_reg[13][29]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][29]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[13][29]~q ),
	.datac(\my_reg[12][29]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux2~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~17 .lut_mask = 16'hAAD8;
defparam \Mux2~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N18
cycloneive_lcell_comb \Mux2~18 (
// Equation(s):
// \Mux2~18_combout  = (dcifimemload_22 & ((\Mux2~17_combout  & ((\my_reg[15][29]~q ))) # (!\Mux2~17_combout  & (\my_reg[14][29]~q )))) # (!dcifimemload_22 & (((\Mux2~17_combout ))))

	.dataa(\my_reg[14][29]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[15][29]~q ),
	.datad(\Mux2~17_combout ),
	.cin(gnd),
	.combout(\Mux2~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~18 .lut_mask = 16'hF388;
defparam \Mux2~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N20
cycloneive_lcell_comb \Mux2~19 (
// Equation(s):
// \Mux2~19_combout  = (\Mux2~16_combout  & (((\Mux2~18_combout )) # (!dcifimemload_24))) # (!\Mux2~16_combout  & (dcifimemload_24 & (\Mux2~11_combout )))

	.dataa(\Mux2~16_combout ),
	.datab(dcifimemload_24),
	.datac(\Mux2~11_combout ),
	.datad(\Mux2~18_combout ),
	.cin(gnd),
	.combout(\Mux2~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~19 .lut_mask = 16'hEA62;
defparam \Mux2~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N21
dffeas \my_reg[27][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][29] .is_wysiwyg = "true";
defparam \my_reg[27][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N19
dffeas \my_reg[31][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][29] .is_wysiwyg = "true";
defparam \my_reg[31][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N17
dffeas \my_reg[19][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][29] .is_wysiwyg = "true";
defparam \my_reg[19][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N16
cycloneive_lcell_comb \Mux2~7 (
// Equation(s):
// \Mux2~7_combout  = (dcifimemload_23 & ((\my_reg[23][29]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[19][29]~q  & !dcifimemload_24))))

	.dataa(\my_reg[23][29]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[19][29]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~7 .lut_mask = 16'hCCB8;
defparam \Mux2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N18
cycloneive_lcell_comb \Mux2~8 (
// Equation(s):
// \Mux2~8_combout  = (dcifimemload_24 & ((\Mux2~7_combout  & ((\my_reg[31][29]~q ))) # (!\Mux2~7_combout  & (\my_reg[27][29]~q )))) # (!dcifimemload_24 & (((\Mux2~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[27][29]~q ),
	.datac(\my_reg[31][29]~q ),
	.datad(\Mux2~7_combout ),
	.cin(gnd),
	.combout(\Mux2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~8 .lut_mask = 16'hF588;
defparam \Mux2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N26
cycloneive_lcell_comb \my_reg[25][29]~feeder (
// Equation(s):
// \my_reg[25][29]~feeder_combout  = \wdat~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat4),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[25][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][29]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[25][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N27
dffeas \my_reg[25][29] (
	.clk(CLK),
	.d(\my_reg[25][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][29] .is_wysiwyg = "true";
defparam \my_reg[25][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N0
cycloneive_lcell_comb \my_reg[21][29]~feeder (
// Equation(s):
// \my_reg[21][29]~feeder_combout  = \wdat~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat4),
	.cin(gnd),
	.combout(\my_reg[21][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][29]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[21][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N1
dffeas \my_reg[21][29] (
	.clk(CLK),
	.d(\my_reg[21][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][29] .is_wysiwyg = "true";
defparam \my_reg[21][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N28
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\my_reg[21][29]~q ))) # (!dcifimemload_23 & (\my_reg[17][29]~q ))))

	.dataa(\my_reg[17][29]~q ),
	.datab(\my_reg[21][29]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hFC0A;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N2
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// \Mux2~1_combout  = (dcifimemload_24 & ((\Mux2~0_combout  & (\my_reg[29][29]~q )) # (!\Mux2~0_combout  & ((\my_reg[25][29]~q ))))) # (!dcifimemload_24 & (((\Mux2~0_combout ))))

	.dataa(\my_reg[29][29]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[25][29]~q ),
	.datad(\Mux2~0_combout ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hBBC0;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N5
dffeas \my_reg[20][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][29] .is_wysiwyg = "true";
defparam \my_reg[20][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N7
dffeas \my_reg[28][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][29] .is_wysiwyg = "true";
defparam \my_reg[28][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N30
cycloneive_lcell_comb \my_reg[24][29]~feeder (
// Equation(s):
// \my_reg[24][29]~feeder_combout  = \wdat~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat4),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[24][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[24][29]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[24][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N31
dffeas \my_reg[24][29] (
	.clk(CLK),
	.d(\my_reg[24][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][29] .is_wysiwyg = "true";
defparam \my_reg[24][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N25
dffeas \my_reg[16][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][29] .is_wysiwyg = "true";
defparam \my_reg[16][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N24
cycloneive_lcell_comb \Mux2~4 (
// Equation(s):
// \Mux2~4_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[24][29]~q )) # (!dcifimemload_24 & ((\my_reg[16][29]~q )))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[24][29]~q ),
	.datac(\my_reg[16][29]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~4 .lut_mask = 16'hEE50;
defparam \Mux2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N6
cycloneive_lcell_comb \Mux2~5 (
// Equation(s):
// \Mux2~5_combout  = (dcifimemload_23 & ((\Mux2~4_combout  & ((\my_reg[28][29]~q ))) # (!\Mux2~4_combout  & (\my_reg[20][29]~q )))) # (!dcifimemload_23 & (((\Mux2~4_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[20][29]~q ),
	.datac(\my_reg[28][29]~q ),
	.datad(\Mux2~4_combout ),
	.cin(gnd),
	.combout(\Mux2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~5 .lut_mask = 16'hF588;
defparam \Mux2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y42_N5
dffeas \my_reg[30][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][29] .is_wysiwyg = "true";
defparam \my_reg[30][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N11
dffeas \my_reg[26][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][29] .is_wysiwyg = "true";
defparam \my_reg[26][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N2
cycloneive_lcell_comb \Mux2~2 (
// Equation(s):
// \Mux2~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\my_reg[26][29]~q ))) # (!dcifimemload_24 & (\my_reg[18][29]~q ))))

	.dataa(\my_reg[18][29]~q ),
	.datab(\my_reg[26][29]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~2 .lut_mask = 16'hFC0A;
defparam \Mux2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N4
cycloneive_lcell_comb \Mux2~3 (
// Equation(s):
// \Mux2~3_combout  = (dcifimemload_23 & ((\Mux2~2_combout  & ((\my_reg[30][29]~q ))) # (!\Mux2~2_combout  & (\my_reg[22][29]~q )))) # (!dcifimemload_23 & (((\Mux2~2_combout ))))

	.dataa(\my_reg[22][29]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[30][29]~q ),
	.datad(\Mux2~2_combout ),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~3 .lut_mask = 16'hF388;
defparam \Mux2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N2
cycloneive_lcell_comb \Mux2~6 (
// Equation(s):
// \Mux2~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux2~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & (\Mux2~5_combout )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux2~5_combout ),
	.datad(\Mux2~3_combout ),
	.cin(gnd),
	.combout(\Mux2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~6 .lut_mask = 16'hBA98;
defparam \Mux2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N8
cycloneive_lcell_comb \Mux2~9 (
// Equation(s):
// \Mux2~9_combout  = (dcifimemload_21 & ((\Mux2~6_combout  & (\Mux2~8_combout )) # (!\Mux2~6_combout  & ((\Mux2~1_combout ))))) # (!dcifimemload_21 & (((\Mux2~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux2~8_combout ),
	.datac(\Mux2~1_combout ),
	.datad(\Mux2~6_combout ),
	.cin(gnd),
	.combout(\Mux2~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~9 .lut_mask = 16'hDDA0;
defparam \Mux2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N14
cycloneive_lcell_comb \Mux34~0 (
// Equation(s):
// \Mux34~0_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][29]~q ))) # (!dcifimemload_16 & (\my_reg[4][29]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[4][29]~q ),
	.datac(\my_reg[5][29]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux34~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~0 .lut_mask = 16'hFA44;
defparam \Mux34~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N24
cycloneive_lcell_comb \Mux34~1 (
// Equation(s):
// \Mux34~1_combout  = (dcifimemload_17 & ((\Mux34~0_combout  & ((\my_reg[7][29]~q ))) # (!\Mux34~0_combout  & (\my_reg[6][29]~q )))) # (!dcifimemload_17 & (\Mux34~0_combout ))

	.dataa(dcifimemload_17),
	.datab(\Mux34~0_combout ),
	.datac(\my_reg[6][29]~q ),
	.datad(\my_reg[7][29]~q ),
	.cin(gnd),
	.combout(\Mux34~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~1 .lut_mask = 16'hEC64;
defparam \Mux34~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N13
dffeas \my_reg[14][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][29] .is_wysiwyg = "true";
defparam \my_reg[14][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N22
cycloneive_lcell_comb \Mux34~7 (
// Equation(s):
// \Mux34~7_combout  = (dcifimemload_16 & (((\my_reg[13][29]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[12][29]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[12][29]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[13][29]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux34~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~7 .lut_mask = 16'hCCE2;
defparam \Mux34~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N12
cycloneive_lcell_comb \Mux34~8 (
// Equation(s):
// \Mux34~8_combout  = (dcifimemload_17 & ((\Mux34~7_combout  & (\my_reg[15][29]~q )) # (!\Mux34~7_combout  & ((\my_reg[14][29]~q ))))) # (!dcifimemload_17 & (((\Mux34~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[15][29]~q ),
	.datac(\my_reg[14][29]~q ),
	.datad(\Mux34~7_combout ),
	.cin(gnd),
	.combout(\Mux34~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~8 .lut_mask = 16'hDDA0;
defparam \Mux34~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N24
cycloneive_lcell_comb \Mux34~2 (
// Equation(s):
// \Mux34~2_combout  = (dcifimemload_17 & (((\my_reg[10][29]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\my_reg[8][29]~q  & ((!dcifimemload_16))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[8][29]~q ),
	.datac(\my_reg[10][29]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux34~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~2 .lut_mask = 16'hAAE4;
defparam \Mux34~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y42_N15
dffeas \my_reg[9][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][29] .is_wysiwyg = "true";
defparam \my_reg[9][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N14
cycloneive_lcell_comb \Mux34~3 (
// Equation(s):
// \Mux34~3_combout  = (\Mux34~2_combout  & ((\my_reg[11][29]~q ) # ((!dcifimemload_16)))) # (!\Mux34~2_combout  & (((\my_reg[9][29]~q  & dcifimemload_16))))

	.dataa(\my_reg[11][29]~q ),
	.datab(\Mux34~2_combout ),
	.datac(\my_reg[9][29]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux34~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~3 .lut_mask = 16'hB8CC;
defparam \Mux34~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N2
cycloneive_lcell_comb \my_reg[1][29]~feeder (
// Equation(s):
// \my_reg[1][29]~feeder_combout  = \wdat~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat4),
	.cin(gnd),
	.combout(\my_reg[1][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[1][29]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[1][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y42_N3
dffeas \my_reg[1][29] (
	.clk(CLK),
	.d(\my_reg[1][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][29] .is_wysiwyg = "true";
defparam \my_reg[1][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N28
cycloneive_lcell_comb \Mux34~4 (
// Equation(s):
// \Mux34~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][29]~q ))) # (!dcifimemload_17 & (\my_reg[1][29]~q ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[1][29]~q ),
	.datac(\my_reg[3][29]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux34~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~4 .lut_mask = 16'hA088;
defparam \Mux34~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N12
cycloneive_lcell_comb \Mux34~5 (
// Equation(s):
// \Mux34~5_combout  = (\Mux34~4_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \my_reg[2][29]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\my_reg[2][29]~q ),
	.datad(\Mux34~4_combout ),
	.cin(gnd),
	.combout(\Mux34~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~5 .lut_mask = 16'hFF40;
defparam \Mux34~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N10
cycloneive_lcell_comb \Mux34~6 (
// Equation(s):
// \Mux34~6_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\Mux34~3_combout )))) # (!dcifimemload_19 & (!dcifimemload_18 & ((\Mux34~5_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux34~3_combout ),
	.datad(\Mux34~5_combout ),
	.cin(gnd),
	.combout(\Mux34~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~6 .lut_mask = 16'hB9A8;
defparam \Mux34~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N2
cycloneive_lcell_comb \Mux34~10 (
// Equation(s):
// \Mux34~10_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[25][29]~q ))) # (!dcifimemload_19 & (\my_reg[17][29]~q ))))

	.dataa(\my_reg[17][29]~q ),
	.datab(\my_reg[25][29]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux34~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~10 .lut_mask = 16'hFC0A;
defparam \Mux34~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N21
dffeas \my_reg[29][29] (
	.clk(CLK),
	.d(wdat4),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][29] .is_wysiwyg = "true";
defparam \my_reg[29][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N20
cycloneive_lcell_comb \Mux34~11 (
// Equation(s):
// \Mux34~11_combout  = (\Mux34~10_combout  & (((\my_reg[29][29]~q ) # (!dcifimemload_18)))) # (!\Mux34~10_combout  & (\my_reg[21][29]~q  & (dcifimemload_18)))

	.dataa(\my_reg[21][29]~q ),
	.datab(\Mux34~10_combout ),
	.datac(dcifimemload_18),
	.datad(\my_reg[29][29]~q ),
	.cin(gnd),
	.combout(\Mux34~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~11 .lut_mask = 16'hEC2C;
defparam \Mux34~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N12
cycloneive_lcell_comb \my_reg[18][29]~feeder (
// Equation(s):
// \my_reg[18][29]~feeder_combout  = \wdat~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat4),
	.cin(gnd),
	.combout(\my_reg[18][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[18][29]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[18][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y42_N13
dffeas \my_reg[18][29] (
	.clk(CLK),
	.d(\my_reg[18][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][29] .is_wysiwyg = "true";
defparam \my_reg[18][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N25
dffeas \my_reg[22][29] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][29] .is_wysiwyg = "true";
defparam \my_reg[22][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N24
cycloneive_lcell_comb \Mux34~12 (
// Equation(s):
// \Mux34~12_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[22][29]~q ))) # (!dcifimemload_18 & (\my_reg[18][29]~q ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[18][29]~q ),
	.datac(\my_reg[22][29]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux34~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~12 .lut_mask = 16'hFA44;
defparam \Mux34~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N10
cycloneive_lcell_comb \Mux34~13 (
// Equation(s):
// \Mux34~13_combout  = (dcifimemload_19 & ((\Mux34~12_combout  & (\my_reg[30][29]~q )) # (!\Mux34~12_combout  & ((\my_reg[26][29]~q ))))) # (!dcifimemload_19 & (((\Mux34~12_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[30][29]~q ),
	.datac(\my_reg[26][29]~q ),
	.datad(\Mux34~12_combout ),
	.cin(gnd),
	.combout(\Mux34~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~13 .lut_mask = 16'hDDA0;
defparam \Mux34~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N4
cycloneive_lcell_comb \Mux34~14 (
// Equation(s):
// \Mux34~14_combout  = (dcifimemload_18 & (((\my_reg[20][29]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[16][29]~q  & ((!dcifimemload_19))))

	.dataa(\my_reg[16][29]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[20][29]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux34~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~14 .lut_mask = 16'hCCE2;
defparam \Mux34~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N24
cycloneive_lcell_comb \Mux34~15 (
// Equation(s):
// \Mux34~15_combout  = (\Mux34~14_combout  & (((\my_reg[28][29]~q ) # (!dcifimemload_19)))) # (!\Mux34~14_combout  & (\my_reg[24][29]~q  & ((dcifimemload_19))))

	.dataa(\my_reg[24][29]~q ),
	.datab(\my_reg[28][29]~q ),
	.datac(\Mux34~14_combout ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux34~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~15 .lut_mask = 16'hCAF0;
defparam \Mux34~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N14
cycloneive_lcell_comb \Mux34~16 (
// Equation(s):
// \Mux34~16_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & (\Mux34~13_combout )) # (!dcifimemload_17 & ((\Mux34~15_combout )))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux34~13_combout ),
	.datad(\Mux34~15_combout ),
	.cin(gnd),
	.combout(\Mux34~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~16 .lut_mask = 16'hD9C8;
defparam \Mux34~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N12
cycloneive_lcell_comb \my_reg[23][29]~feeder (
// Equation(s):
// \my_reg[23][29]~feeder_combout  = \wdat~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat4),
	.cin(gnd),
	.combout(\my_reg[23][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[23][29]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[23][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N13
dffeas \my_reg[23][29] (
	.clk(CLK),
	.d(\my_reg[23][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][29] .is_wysiwyg = "true";
defparam \my_reg[23][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N20
cycloneive_lcell_comb \Mux34~17 (
// Equation(s):
// \Mux34~17_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\my_reg[27][29]~q )))) # (!dcifimemload_19 & (!dcifimemload_18 & ((\my_reg[19][29]~q ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\my_reg[27][29]~q ),
	.datad(\my_reg[19][29]~q ),
	.cin(gnd),
	.combout(\Mux34~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~17 .lut_mask = 16'hB9A8;
defparam \Mux34~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N6
cycloneive_lcell_comb \Mux34~18 (
// Equation(s):
// \Mux34~18_combout  = (dcifimemload_18 & ((\Mux34~17_combout  & ((\my_reg[31][29]~q ))) # (!\Mux34~17_combout  & (\my_reg[23][29]~q )))) # (!dcifimemload_18 & (((\Mux34~17_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[23][29]~q ),
	.datac(\my_reg[31][29]~q ),
	.datad(\Mux34~17_combout ),
	.cin(gnd),
	.combout(\Mux34~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~18 .lut_mask = 16'hF588;
defparam \Mux34~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N9
dffeas \my_reg[2][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][28] .is_wysiwyg = "true";
defparam \my_reg[2][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N19
dffeas \my_reg[1][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][28] .is_wysiwyg = "true";
defparam \my_reg[1][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y42_N9
dffeas \my_reg[3][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][28] .is_wysiwyg = "true";
defparam \my_reg[3][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N18
cycloneive_lcell_comb \Mux3~14 (
// Equation(s):
// \Mux3~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][28]~q ))) # (!dcifimemload_22 & (\my_reg[1][28]~q ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\my_reg[1][28]~q ),
	.datad(\my_reg[3][28]~q ),
	.cin(gnd),
	.combout(\Mux3~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~14 .lut_mask = 16'hC840;
defparam \Mux3~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N8
cycloneive_lcell_comb \Mux3~15 (
// Equation(s):
// \Mux3~15_combout  = (\Mux3~14_combout ) # ((dcifimemload_22 & (!dcifimemload_21 & \my_reg[2][28]~q )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\my_reg[2][28]~q ),
	.datad(\Mux3~14_combout ),
	.cin(gnd),
	.combout(\Mux3~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~15 .lut_mask = 16'hFF20;
defparam \Mux3~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y42_N27
dffeas \my_reg[9][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][28] .is_wysiwyg = "true";
defparam \my_reg[9][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N3
dffeas \my_reg[11][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][28] .is_wysiwyg = "true";
defparam \my_reg[11][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y42_N29
dffeas \my_reg[10][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][28] .is_wysiwyg = "true";
defparam \my_reg[10][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N17
dffeas \my_reg[8][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][28] .is_wysiwyg = "true";
defparam \my_reg[8][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N16
cycloneive_lcell_comb \Mux3~12 (
// Equation(s):
// \Mux3~12_combout  = (dcifimemload_22 & ((\my_reg[10][28]~q ) # ((dcifimemload_21)))) # (!dcifimemload_22 & (((\my_reg[8][28]~q  & !dcifimemload_21))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[10][28]~q ),
	.datac(\my_reg[8][28]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux3~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~12 .lut_mask = 16'hAAD8;
defparam \Mux3~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N2
cycloneive_lcell_comb \Mux3~13 (
// Equation(s):
// \Mux3~13_combout  = (dcifimemload_21 & ((\Mux3~12_combout  & ((\my_reg[11][28]~q ))) # (!\Mux3~12_combout  & (\my_reg[9][28]~q )))) # (!dcifimemload_21 & (((\Mux3~12_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][28]~q ),
	.datac(\my_reg[11][28]~q ),
	.datad(\Mux3~12_combout ),
	.cin(gnd),
	.combout(\Mux3~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~13 .lut_mask = 16'hF588;
defparam \Mux3~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N10
cycloneive_lcell_comb \Mux3~16 (
// Equation(s):
// \Mux3~16_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\Mux3~13_combout ))) # (!dcifimemload_24 & (\Mux3~15_combout ))))

	.dataa(dcifimemload_23),
	.datab(\Mux3~15_combout ),
	.datac(dcifimemload_24),
	.datad(\Mux3~13_combout ),
	.cin(gnd),
	.combout(\Mux3~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~16 .lut_mask = 16'hF4A4;
defparam \Mux3~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N15
dffeas \my_reg[15][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][28] .is_wysiwyg = "true";
defparam \my_reg[15][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y41_N29
dffeas \my_reg[14][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][28] .is_wysiwyg = "true";
defparam \my_reg[14][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N14
cycloneive_lcell_comb \Mux3~18 (
// Equation(s):
// \Mux3~18_combout  = (\Mux3~17_combout  & (((\my_reg[15][28]~q )) # (!dcifimemload_22))) # (!\Mux3~17_combout  & (dcifimemload_22 & ((\my_reg[14][28]~q ))))

	.dataa(\Mux3~17_combout ),
	.datab(dcifimemload_22),
	.datac(\my_reg[15][28]~q ),
	.datad(\my_reg[14][28]~q ),
	.cin(gnd),
	.combout(\Mux3~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~18 .lut_mask = 16'hE6A2;
defparam \Mux3~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N13
dffeas \my_reg[6][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][28] .is_wysiwyg = "true";
defparam \my_reg[6][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N15
dffeas \my_reg[7][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][28] .is_wysiwyg = "true";
defparam \my_reg[7][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y42_N11
dffeas \my_reg[5][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][28] .is_wysiwyg = "true";
defparam \my_reg[5][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N29
dffeas \my_reg[4][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][28] .is_wysiwyg = "true";
defparam \my_reg[4][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N28
cycloneive_lcell_comb \Mux3~10 (
// Equation(s):
// \Mux3~10_combout  = (dcifimemload_21 & ((\my_reg[5][28]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[4][28]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[5][28]~q ),
	.datac(\my_reg[4][28]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux3~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~10 .lut_mask = 16'hAAD8;
defparam \Mux3~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N14
cycloneive_lcell_comb \Mux3~11 (
// Equation(s):
// \Mux3~11_combout  = (dcifimemload_22 & ((\Mux3~10_combout  & ((\my_reg[7][28]~q ))) # (!\Mux3~10_combout  & (\my_reg[6][28]~q )))) # (!dcifimemload_22 & (((\Mux3~10_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[6][28]~q ),
	.datac(\my_reg[7][28]~q ),
	.datad(\Mux3~10_combout ),
	.cin(gnd),
	.combout(\Mux3~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~11 .lut_mask = 16'hF588;
defparam \Mux3~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N24
cycloneive_lcell_comb \Mux3~19 (
// Equation(s):
// \Mux3~19_combout  = (\Mux3~16_combout  & (((\Mux3~18_combout )) # (!dcifimemload_23))) # (!\Mux3~16_combout  & (dcifimemload_23 & ((\Mux3~11_combout ))))

	.dataa(\Mux3~16_combout ),
	.datab(dcifimemload_23),
	.datac(\Mux3~18_combout ),
	.datad(\Mux3~11_combout ),
	.cin(gnd),
	.combout(\Mux3~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~19 .lut_mask = 16'hE6A2;
defparam \Mux3~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N5
dffeas \my_reg[19][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][28] .is_wysiwyg = "true";
defparam \my_reg[19][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N4
cycloneive_lcell_comb \Mux3~7 (
// Equation(s):
// \Mux3~7_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[27][28]~q )) # (!dcifimemload_24 & ((\my_reg[19][28]~q )))))

	.dataa(\my_reg[27][28]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[19][28]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~7 .lut_mask = 16'hEE30;
defparam \Mux3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N31
dffeas \my_reg[31][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][28] .is_wysiwyg = "true";
defparam \my_reg[31][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N30
cycloneive_lcell_comb \Mux3~8 (
// Equation(s):
// \Mux3~8_combout  = (\Mux3~7_combout  & (((\my_reg[31][28]~q ) # (!dcifimemload_23)))) # (!\Mux3~7_combout  & (\my_reg[23][28]~q  & ((dcifimemload_23))))

	.dataa(\my_reg[23][28]~q ),
	.datab(\Mux3~7_combout ),
	.datac(\my_reg[31][28]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux3~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~8 .lut_mask = 16'hE2CC;
defparam \Mux3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N1
dffeas \my_reg[26][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][28] .is_wysiwyg = "true";
defparam \my_reg[26][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y42_N23
dffeas \my_reg[30][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][28] .is_wysiwyg = "true";
defparam \my_reg[30][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N24
cycloneive_lcell_comb \my_reg[18][28]~feeder (
// Equation(s):
// \my_reg[18][28]~feeder_combout  = \wdat~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat5),
	.cin(gnd),
	.combout(\my_reg[18][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[18][28]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[18][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N25
dffeas \my_reg[18][28] (
	.clk(CLK),
	.d(\my_reg[18][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][28] .is_wysiwyg = "true";
defparam \my_reg[18][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N23
dffeas \my_reg[22][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][28] .is_wysiwyg = "true";
defparam \my_reg[22][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N10
cycloneive_lcell_comb \Mux3~2 (
// Equation(s):
// \Mux3~2_combout  = (dcifimemload_23 & (((\my_reg[22][28]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\my_reg[18][28]~q  & ((!dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[18][28]~q ),
	.datac(\my_reg[22][28]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~2 .lut_mask = 16'hAAE4;
defparam \Mux3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N22
cycloneive_lcell_comb \Mux3~3 (
// Equation(s):
// \Mux3~3_combout  = (dcifimemload_24 & ((\Mux3~2_combout  & ((\my_reg[30][28]~q ))) # (!\Mux3~2_combout  & (\my_reg[26][28]~q )))) # (!dcifimemload_24 & (((\Mux3~2_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[26][28]~q ),
	.datac(\my_reg[30][28]~q ),
	.datad(\Mux3~2_combout ),
	.cin(gnd),
	.combout(\Mux3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~3 .lut_mask = 16'hF588;
defparam \Mux3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y40_N15
dffeas \my_reg[24][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][28] .is_wysiwyg = "true";
defparam \my_reg[24][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N27
dffeas \my_reg[28][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][28] .is_wysiwyg = "true";
defparam \my_reg[28][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y40_N1
dffeas \my_reg[20][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][28] .is_wysiwyg = "true";
defparam \my_reg[20][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N1
dffeas \my_reg[16][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][28] .is_wysiwyg = "true";
defparam \my_reg[16][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N0
cycloneive_lcell_comb \Mux3~4 (
// Equation(s):
// \Mux3~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[20][28]~q )) # (!dcifimemload_23 & ((\my_reg[16][28]~q )))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[20][28]~q ),
	.datac(\my_reg[16][28]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~4 .lut_mask = 16'hEE50;
defparam \Mux3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N26
cycloneive_lcell_comb \Mux3~5 (
// Equation(s):
// \Mux3~5_combout  = (dcifimemload_24 & ((\Mux3~4_combout  & ((\my_reg[28][28]~q ))) # (!\Mux3~4_combout  & (\my_reg[24][28]~q )))) # (!dcifimemload_24 & (((\Mux3~4_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[24][28]~q ),
	.datac(\my_reg[28][28]~q ),
	.datad(\Mux3~4_combout ),
	.cin(gnd),
	.combout(\Mux3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~5 .lut_mask = 16'hF588;
defparam \Mux3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N22
cycloneive_lcell_comb \Mux3~6 (
// Equation(s):
// \Mux3~6_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\Mux3~3_combout )) # (!dcifimemload_22 & ((\Mux3~5_combout )))))

	.dataa(dcifimemload_21),
	.datab(\Mux3~3_combout ),
	.datac(dcifimemload_22),
	.datad(\Mux3~5_combout ),
	.cin(gnd),
	.combout(\Mux3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~6 .lut_mask = 16'hE5E0;
defparam \Mux3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N7
dffeas \my_reg[29][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][28] .is_wysiwyg = "true";
defparam \my_reg[29][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N1
dffeas \my_reg[17][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][28] .is_wysiwyg = "true";
defparam \my_reg[17][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N0
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[25][28]~q )) # (!dcifimemload_24 & ((\my_reg[17][28]~q )))))

	.dataa(\my_reg[25][28]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[17][28]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hEE30;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N6
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (dcifimemload_23 & ((\Mux3~0_combout  & ((\my_reg[29][28]~q ))) # (!\Mux3~0_combout  & (\my_reg[21][28]~q )))) # (!dcifimemload_23 & (((\Mux3~0_combout ))))

	.dataa(\my_reg[21][28]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[29][28]~q ),
	.datad(\Mux3~0_combout ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hF388;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N16
cycloneive_lcell_comb \Mux3~9 (
// Equation(s):
// \Mux3~9_combout  = (dcifimemload_21 & ((\Mux3~6_combout  & (\Mux3~8_combout )) # (!\Mux3~6_combout  & ((\Mux3~1_combout ))))) # (!dcifimemload_21 & (((\Mux3~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux3~8_combout ),
	.datac(\Mux3~6_combout ),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\Mux3~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~9 .lut_mask = 16'hDAD0;
defparam \Mux3~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N29
dffeas \my_reg[13][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][28] .is_wysiwyg = "true";
defparam \my_reg[13][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N28
cycloneive_lcell_comb \Mux35~7 (
// Equation(s):
// \Mux35~7_combout  = (dcifimemload_16 & (((\my_reg[13][28]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[12][28]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[12][28]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[13][28]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux35~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~7 .lut_mask = 16'hCCE2;
defparam \Mux35~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N28
cycloneive_lcell_comb \Mux35~8 (
// Equation(s):
// \Mux35~8_combout  = (dcifimemload_17 & ((\Mux35~7_combout  & (\my_reg[15][28]~q )) # (!\Mux35~7_combout  & ((\my_reg[14][28]~q ))))) # (!dcifimemload_17 & (((\Mux35~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[15][28]~q ),
	.datac(\my_reg[14][28]~q ),
	.datad(\Mux35~7_combout ),
	.cin(gnd),
	.combout(\Mux35~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~8 .lut_mask = 16'hDDA0;
defparam \Mux35~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N8
cycloneive_lcell_comb \Mux35~4 (
// Equation(s):
// \Mux35~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][28]~q ))) # (!dcifimemload_17 & (\my_reg[1][28]~q ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[1][28]~q ),
	.datac(\my_reg[3][28]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux35~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~4 .lut_mask = 16'hA088;
defparam \Mux35~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N22
cycloneive_lcell_comb \Mux35~5 (
// Equation(s):
// \Mux35~5_combout  = (\Mux35~4_combout ) # ((!dcifimemload_16 & (\my_reg[2][28]~q  & dcifimemload_17)))

	.dataa(dcifimemload_16),
	.datab(\my_reg[2][28]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux35~4_combout ),
	.cin(gnd),
	.combout(\Mux35~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~5 .lut_mask = 16'hFF40;
defparam \Mux35~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N10
cycloneive_lcell_comb \Mux35~2 (
// Equation(s):
// \Mux35~2_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][28]~q ))) # (!dcifimemload_16 & (\my_reg[4][28]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[4][28]~q ),
	.datac(\my_reg[5][28]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux35~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~2 .lut_mask = 16'hFA44;
defparam \Mux35~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N12
cycloneive_lcell_comb \Mux35~3 (
// Equation(s):
// \Mux35~3_combout  = (dcifimemload_17 & ((\Mux35~2_combout  & (\my_reg[7][28]~q )) # (!\Mux35~2_combout  & ((\my_reg[6][28]~q ))))) # (!dcifimemload_17 & (((\Mux35~2_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[7][28]~q ),
	.datac(\my_reg[6][28]~q ),
	.datad(\Mux35~2_combout ),
	.cin(gnd),
	.combout(\Mux35~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~3 .lut_mask = 16'hDDA0;
defparam \Mux35~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N8
cycloneive_lcell_comb \Mux35~6 (
// Equation(s):
// \Mux35~6_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & ((\Mux35~3_combout ))) # (!dcifimemload_18 & (\Mux35~5_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux35~5_combout ),
	.datad(\Mux35~3_combout ),
	.cin(gnd),
	.combout(\Mux35~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~6 .lut_mask = 16'hDC98;
defparam \Mux35~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N28
cycloneive_lcell_comb \Mux35~0 (
// Equation(s):
// \Mux35~0_combout  = (dcifimemload_17 & (((\my_reg[10][28]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\my_reg[8][28]~q  & ((!dcifimemload_16))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[8][28]~q ),
	.datac(\my_reg[10][28]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux35~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~0 .lut_mask = 16'hAAE4;
defparam \Mux35~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N26
cycloneive_lcell_comb \Mux35~1 (
// Equation(s):
// \Mux35~1_combout  = (\Mux35~0_combout  & ((\my_reg[11][28]~q ) # ((!dcifimemload_16)))) # (!\Mux35~0_combout  & (((\my_reg[9][28]~q  & dcifimemload_16))))

	.dataa(\my_reg[11][28]~q ),
	.datab(\Mux35~0_combout ),
	.datac(\my_reg[9][28]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux35~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~1 .lut_mask = 16'hB8CC;
defparam \Mux35~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N2
cycloneive_lcell_comb \my_reg[25][28]~feeder (
// Equation(s):
// \my_reg[25][28]~feeder_combout  = \wdat~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat5),
	.cin(gnd),
	.combout(\my_reg[25][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][28]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[25][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N3
dffeas \my_reg[25][28] (
	.clk(CLK),
	.d(\my_reg[25][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][28] .is_wysiwyg = "true";
defparam \my_reg[25][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N6
cycloneive_lcell_comb \Mux35~10 (
// Equation(s):
// \Mux35~10_combout  = (dcifimemload_18 & ((\my_reg[21][28]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((!dcifimemload_19 & \my_reg[17][28]~q ))))

	.dataa(\my_reg[21][28]~q ),
	.datab(dcifimemload_18),
	.datac(dcifimemload_19),
	.datad(\my_reg[17][28]~q ),
	.cin(gnd),
	.combout(\Mux35~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~10 .lut_mask = 16'hCBC8;
defparam \Mux35~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N12
cycloneive_lcell_comb \Mux35~11 (
// Equation(s):
// \Mux35~11_combout  = (dcifimemload_19 & ((\Mux35~10_combout  & ((\my_reg[29][28]~q ))) # (!\Mux35~10_combout  & (\my_reg[25][28]~q )))) # (!dcifimemload_19 & (((\Mux35~10_combout ))))

	.dataa(\my_reg[25][28]~q ),
	.datab(\my_reg[29][28]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux35~10_combout ),
	.cin(gnd),
	.combout(\Mux35~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~11 .lut_mask = 16'hCFA0;
defparam \Mux35~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N25
dffeas \my_reg[27][28] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][28] .is_wysiwyg = "true";
defparam \my_reg[27][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N10
cycloneive_lcell_comb \my_reg[23][28]~feeder (
// Equation(s):
// \my_reg[23][28]~feeder_combout  = \wdat~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat5),
	.cin(gnd),
	.combout(\my_reg[23][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[23][28]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[23][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N11
dffeas \my_reg[23][28] (
	.clk(CLK),
	.d(\my_reg[23][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][28] .is_wysiwyg = "true";
defparam \my_reg[23][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N10
cycloneive_lcell_comb \Mux35~17 (
// Equation(s):
// \Mux35~17_combout  = (dcifimemload_18 & (((dcifimemload_19) # (\my_reg[23][28]~q )))) # (!dcifimemload_18 & (\my_reg[19][28]~q  & (!dcifimemload_19)))

	.dataa(\my_reg[19][28]~q ),
	.datab(dcifimemload_18),
	.datac(dcifimemload_19),
	.datad(\my_reg[23][28]~q ),
	.cin(gnd),
	.combout(\Mux35~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~17 .lut_mask = 16'hCEC2;
defparam \Mux35~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N24
cycloneive_lcell_comb \Mux35~18 (
// Equation(s):
// \Mux35~18_combout  = (dcifimemload_19 & ((\Mux35~17_combout  & (\my_reg[31][28]~q )) # (!\Mux35~17_combout  & ((\my_reg[27][28]~q ))))) # (!dcifimemload_19 & (((\Mux35~17_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[31][28]~q ),
	.datac(\my_reg[27][28]~q ),
	.datad(\Mux35~17_combout ),
	.cin(gnd),
	.combout(\Mux35~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~18 .lut_mask = 16'hDDA0;
defparam \Mux35~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N14
cycloneive_lcell_comb \Mux35~14 (
// Equation(s):
// \Mux35~14_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & (\my_reg[24][28]~q )) # (!dcifimemload_19 & ((\my_reg[16][28]~q )))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\my_reg[24][28]~q ),
	.datad(\my_reg[16][28]~q ),
	.cin(gnd),
	.combout(\Mux35~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~14 .lut_mask = 16'hD9C8;
defparam \Mux35~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N0
cycloneive_lcell_comb \Mux35~15 (
// Equation(s):
// \Mux35~15_combout  = (dcifimemload_18 & ((\Mux35~14_combout  & (\my_reg[28][28]~q )) # (!\Mux35~14_combout  & ((\my_reg[20][28]~q ))))) # (!dcifimemload_18 & (((\Mux35~14_combout ))))

	.dataa(\my_reg[28][28]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[20][28]~q ),
	.datad(\Mux35~14_combout ),
	.cin(gnd),
	.combout(\Mux35~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~15 .lut_mask = 16'hBBC0;
defparam \Mux35~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N0
cycloneive_lcell_comb \Mux35~12 (
// Equation(s):
// \Mux35~12_combout  = (dcifimemload_19 & (((\my_reg[26][28]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[18][28]~q  & ((!dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[18][28]~q ),
	.datac(\my_reg[26][28]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux35~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~12 .lut_mask = 16'hAAE4;
defparam \Mux35~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N22
cycloneive_lcell_comb \Mux35~13 (
// Equation(s):
// \Mux35~13_combout  = (dcifimemload_18 & ((\Mux35~12_combout  & (\my_reg[30][28]~q )) # (!\Mux35~12_combout  & ((\my_reg[22][28]~q ))))) # (!dcifimemload_18 & (((\Mux35~12_combout ))))

	.dataa(\my_reg[30][28]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[22][28]~q ),
	.datad(\Mux35~12_combout ),
	.cin(gnd),
	.combout(\Mux35~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~13 .lut_mask = 16'hBBC0;
defparam \Mux35~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N26
cycloneive_lcell_comb \Mux35~16 (
// Equation(s):
// \Mux35~16_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux35~13_combout ))) # (!dcifimemload_17 & (\Mux35~15_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux35~15_combout ),
	.datac(dcifimemload_17),
	.datad(\Mux35~13_combout ),
	.cin(gnd),
	.combout(\Mux35~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~16 .lut_mask = 16'hF4A4;
defparam \Mux35~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y42_N13
dffeas \my_reg[25][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][27] .is_wysiwyg = "true";
defparam \my_reg[25][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N25
dffeas \my_reg[29][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][27] .is_wysiwyg = "true";
defparam \my_reg[29][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N11
dffeas \my_reg[17][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][27] .is_wysiwyg = "true";
defparam \my_reg[17][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N10
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (dcifimemload_23 & ((\my_reg[21][27]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[17][27]~q  & !dcifimemload_24))))

	.dataa(\my_reg[21][27]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[17][27]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hCCB8;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N24
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// \Mux4~1_combout  = (dcifimemload_24 & ((\Mux4~0_combout  & ((\my_reg[29][27]~q ))) # (!\Mux4~0_combout  & (\my_reg[25][27]~q )))) # (!dcifimemload_24 & (((\Mux4~0_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[25][27]~q ),
	.datac(\my_reg[29][27]~q ),
	.datad(\Mux4~0_combout ),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hF588;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N24
cycloneive_lcell_comb \my_reg[22][27]~feeder (
// Equation(s):
// \my_reg[22][27]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat6),
	.cin(gnd),
	.combout(\my_reg[22][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[22][27]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[22][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y43_N25
dffeas \my_reg[22][27] (
	.clk(CLK),
	.d(\my_reg[22][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][27] .is_wysiwyg = "true";
defparam \my_reg[22][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N20
cycloneive_lcell_comb \my_reg[26][27]~feeder (
// Equation(s):
// \my_reg[26][27]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat6),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[26][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[26][27]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[26][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N21
dffeas \my_reg[26][27] (
	.clk(CLK),
	.d(\my_reg[26][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][27] .is_wysiwyg = "true";
defparam \my_reg[26][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N2
cycloneive_lcell_comb \my_reg[18][27]~feeder (
// Equation(s):
// \my_reg[18][27]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat6),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[18][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[18][27]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[18][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N3
dffeas \my_reg[18][27] (
	.clk(CLK),
	.d(\my_reg[18][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][27] .is_wysiwyg = "true";
defparam \my_reg[18][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N28
cycloneive_lcell_comb \Mux4~2 (
// Equation(s):
// \Mux4~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[26][27]~q )) # (!dcifimemload_24 & ((\my_reg[18][27]~q )))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[26][27]~q ),
	.datac(\my_reg[18][27]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~2 .lut_mask = 16'hEE50;
defparam \Mux4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N14
cycloneive_lcell_comb \Mux4~3 (
// Equation(s):
// \Mux4~3_combout  = (\Mux4~2_combout  & ((\my_reg[30][27]~q ) # ((!dcifimemload_23)))) # (!\Mux4~2_combout  & (((\my_reg[22][27]~q  & dcifimemload_23))))

	.dataa(\my_reg[30][27]~q ),
	.datab(\my_reg[22][27]~q ),
	.datac(\Mux4~2_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~3 .lut_mask = 16'hACF0;
defparam \Mux4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N18
cycloneive_lcell_comb \my_reg[28][27]~feeder (
// Equation(s):
// \my_reg[28][27]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat6),
	.cin(gnd),
	.combout(\my_reg[28][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[28][27]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[28][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y43_N19
dffeas \my_reg[28][27] (
	.clk(CLK),
	.d(\my_reg[28][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][27] .is_wysiwyg = "true";
defparam \my_reg[28][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N4
cycloneive_lcell_comb \my_reg[16][27]~feeder (
// Equation(s):
// \my_reg[16][27]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat6),
	.cin(gnd),
	.combout(\my_reg[16][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[16][27]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[16][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N5
dffeas \my_reg[16][27] (
	.clk(CLK),
	.d(\my_reg[16][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][27] .is_wysiwyg = "true";
defparam \my_reg[16][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N4
cycloneive_lcell_comb \Mux4~4 (
// Equation(s):
// \Mux4~4_combout  = (dcifimemload_24 & ((\my_reg[24][27]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\my_reg[16][27]~q  & !dcifimemload_23))))

	.dataa(\my_reg[24][27]~q ),
	.datab(\my_reg[16][27]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~4 .lut_mask = 16'hF0AC;
defparam \Mux4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N12
cycloneive_lcell_comb \Mux4~5 (
// Equation(s):
// \Mux4~5_combout  = (\Mux4~4_combout  & (((\my_reg[28][27]~q ) # (!dcifimemload_23)))) # (!\Mux4~4_combout  & (\my_reg[20][27]~q  & ((dcifimemload_23))))

	.dataa(\my_reg[20][27]~q ),
	.datab(\my_reg[28][27]~q ),
	.datac(\Mux4~4_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~5 .lut_mask = 16'hCAF0;
defparam \Mux4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N26
cycloneive_lcell_comb \Mux4~6 (
// Equation(s):
// \Mux4~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux4~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\Mux4~5_combout ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux4~3_combout ),
	.datad(\Mux4~5_combout ),
	.cin(gnd),
	.combout(\Mux4~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~6 .lut_mask = 16'hB9A8;
defparam \Mux4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N25
dffeas \my_reg[27][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][27] .is_wysiwyg = "true";
defparam \my_reg[27][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N3
dffeas \my_reg[31][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][27] .is_wysiwyg = "true";
defparam \my_reg[31][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N21
dffeas \my_reg[19][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][27] .is_wysiwyg = "true";
defparam \my_reg[19][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N20
cycloneive_lcell_comb \Mux4~7 (
// Equation(s):
// \Mux4~7_combout  = (dcifimemload_23 & ((\my_reg[23][27]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[19][27]~q  & !dcifimemload_24))))

	.dataa(\my_reg[23][27]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[19][27]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux4~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~7 .lut_mask = 16'hCCB8;
defparam \Mux4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N2
cycloneive_lcell_comb \Mux4~8 (
// Equation(s):
// \Mux4~8_combout  = (dcifimemload_24 & ((\Mux4~7_combout  & ((\my_reg[31][27]~q ))) # (!\Mux4~7_combout  & (\my_reg[27][27]~q )))) # (!dcifimemload_24 & (((\Mux4~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[27][27]~q ),
	.datac(\my_reg[31][27]~q ),
	.datad(\Mux4~7_combout ),
	.cin(gnd),
	.combout(\Mux4~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~8 .lut_mask = 16'hF588;
defparam \Mux4~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N12
cycloneive_lcell_comb \Mux4~9 (
// Equation(s):
// \Mux4~9_combout  = (dcifimemload_21 & ((\Mux4~6_combout  & ((\Mux4~8_combout ))) # (!\Mux4~6_combout  & (\Mux4~1_combout )))) # (!dcifimemload_21 & (((\Mux4~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux4~1_combout ),
	.datac(\Mux4~6_combout ),
	.datad(\Mux4~8_combout ),
	.cin(gnd),
	.combout(\Mux4~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~9 .lut_mask = 16'hF858;
defparam \Mux4~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N11
dffeas \my_reg[15][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][27] .is_wysiwyg = "true";
defparam \my_reg[15][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N2
cycloneive_lcell_comb \my_reg[13][27]~feeder (
// Equation(s):
// \my_reg[13][27]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat6),
	.cin(gnd),
	.combout(\my_reg[13][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[13][27]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[13][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N3
dffeas \my_reg[13][27] (
	.clk(CLK),
	.d(\my_reg[13][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][27] .is_wysiwyg = "true";
defparam \my_reg[13][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N29
dffeas \my_reg[12][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][27] .is_wysiwyg = "true";
defparam \my_reg[12][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N28
cycloneive_lcell_comb \Mux4~17 (
// Equation(s):
// \Mux4~17_combout  = (dcifimemload_21 & ((\my_reg[13][27]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][27]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[13][27]~q ),
	.datac(\my_reg[12][27]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux4~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~17 .lut_mask = 16'hAAD8;
defparam \Mux4~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N10
cycloneive_lcell_comb \Mux4~18 (
// Equation(s):
// \Mux4~18_combout  = (dcifimemload_22 & ((\Mux4~17_combout  & ((\my_reg[15][27]~q ))) # (!\Mux4~17_combout  & (\my_reg[14][27]~q )))) # (!dcifimemload_22 & (((\Mux4~17_combout ))))

	.dataa(\my_reg[14][27]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[15][27]~q ),
	.datad(\Mux4~17_combout ),
	.cin(gnd),
	.combout(\Mux4~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~18 .lut_mask = 16'hF388;
defparam \Mux4~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N2
cycloneive_lcell_comb \my_reg[9][27]~feeder (
// Equation(s):
// \my_reg[9][27]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat6),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[9][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[9][27]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[9][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N3
dffeas \my_reg[9][27] (
	.clk(CLK),
	.d(\my_reg[9][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][27] .is_wysiwyg = "true";
defparam \my_reg[9][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N28
cycloneive_lcell_comb \my_reg[10][27]~feeder (
// Equation(s):
// \my_reg[10][27]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat6),
	.cin(gnd),
	.combout(\my_reg[10][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[10][27]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[10][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y38_N29
dffeas \my_reg[10][27] (
	.clk(CLK),
	.d(\my_reg[10][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][27] .is_wysiwyg = "true";
defparam \my_reg[10][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N26
cycloneive_lcell_comb \Mux4~10 (
// Equation(s):
// \Mux4~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[10][27]~q ))) # (!dcifimemload_22 & (\my_reg[8][27]~q ))))

	.dataa(\my_reg[8][27]~q ),
	.datab(\my_reg[10][27]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux4~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~10 .lut_mask = 16'hFC0A;
defparam \Mux4~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N16
cycloneive_lcell_comb \Mux4~11 (
// Equation(s):
// \Mux4~11_combout  = (dcifimemload_21 & ((\Mux4~10_combout  & (\my_reg[11][27]~q )) # (!\Mux4~10_combout  & ((\my_reg[9][27]~q ))))) # (!dcifimemload_21 & (((\Mux4~10_combout ))))

	.dataa(\my_reg[11][27]~q ),
	.datab(\my_reg[9][27]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux4~10_combout ),
	.cin(gnd),
	.combout(\Mux4~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~11 .lut_mask = 16'hAFC0;
defparam \Mux4~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N12
cycloneive_lcell_comb \my_reg[7][27]~feeder (
// Equation(s):
// \my_reg[7][27]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat6),
	.cin(gnd),
	.combout(\my_reg[7][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[7][27]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[7][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y43_N13
dffeas \my_reg[7][27] (
	.clk(CLK),
	.d(\my_reg[7][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][27] .is_wysiwyg = "true";
defparam \my_reg[7][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N24
cycloneive_lcell_comb \my_reg[6][27]~feeder (
// Equation(s):
// \my_reg[6][27]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat6),
	.cin(gnd),
	.combout(\my_reg[6][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[6][27]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[6][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y32_N25
dffeas \my_reg[6][27] (
	.clk(CLK),
	.d(\my_reg[6][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][27] .is_wysiwyg = "true";
defparam \my_reg[6][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N4
cycloneive_lcell_comb \my_reg[4][27]~feeder (
// Equation(s):
// \my_reg[4][27]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat6),
	.cin(gnd),
	.combout(\my_reg[4][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[4][27]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[4][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y43_N5
dffeas \my_reg[4][27] (
	.clk(CLK),
	.d(\my_reg[4][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][27] .is_wysiwyg = "true";
defparam \my_reg[4][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N18
cycloneive_lcell_comb \Mux4~12 (
// Equation(s):
// \Mux4~12_combout  = (dcifimemload_21 & ((\my_reg[5][27]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[4][27]~q  & !dcifimemload_22))))

	.dataa(\my_reg[5][27]~q ),
	.datab(\my_reg[4][27]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux4~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~12 .lut_mask = 16'hF0AC;
defparam \Mux4~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N26
cycloneive_lcell_comb \Mux4~13 (
// Equation(s):
// \Mux4~13_combout  = (dcifimemload_22 & ((\Mux4~12_combout  & (\my_reg[7][27]~q )) # (!\Mux4~12_combout  & ((\my_reg[6][27]~q ))))) # (!dcifimemload_22 & (((\Mux4~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[7][27]~q ),
	.datac(\my_reg[6][27]~q ),
	.datad(\Mux4~12_combout ),
	.cin(gnd),
	.combout(\Mux4~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~13 .lut_mask = 16'hDDA0;
defparam \Mux4~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y43_N25
dffeas \my_reg[2][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][27] .is_wysiwyg = "true";
defparam \my_reg[2][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y42_N17
dffeas \my_reg[1][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][27] .is_wysiwyg = "true";
defparam \my_reg[1][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N16
cycloneive_lcell_comb \Mux4~14 (
// Equation(s):
// \Mux4~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\my_reg[3][27]~q )) # (!dcifimemload_22 & ((\my_reg[1][27]~q )))))

	.dataa(\my_reg[3][27]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[1][27]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux4~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~14 .lut_mask = 16'hB800;
defparam \Mux4~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N24
cycloneive_lcell_comb \Mux4~15 (
// Equation(s):
// \Mux4~15_combout  = (\Mux4~14_combout ) # ((!dcifimemload_21 & (dcifimemload_22 & \my_reg[2][27]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\my_reg[2][27]~q ),
	.datad(\Mux4~14_combout ),
	.cin(gnd),
	.combout(\Mux4~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~15 .lut_mask = 16'hFF40;
defparam \Mux4~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N20
cycloneive_lcell_comb \Mux4~16 (
// Equation(s):
// \Mux4~16_combout  = (dcifimemload_23 & ((dcifimemload_24) # ((\Mux4~13_combout )))) # (!dcifimemload_23 & (!dcifimemload_24 & ((\Mux4~15_combout ))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux4~13_combout ),
	.datad(\Mux4~15_combout ),
	.cin(gnd),
	.combout(\Mux4~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~16 .lut_mask = 16'hB9A8;
defparam \Mux4~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N14
cycloneive_lcell_comb \Mux4~19 (
// Equation(s):
// \Mux4~19_combout  = (dcifimemload_24 & ((\Mux4~16_combout  & (\Mux4~18_combout )) # (!\Mux4~16_combout  & ((\Mux4~11_combout ))))) # (!dcifimemload_24 & (((\Mux4~16_combout ))))

	.dataa(\Mux4~18_combout ),
	.datab(dcifimemload_24),
	.datac(\Mux4~11_combout ),
	.datad(\Mux4~16_combout ),
	.cin(gnd),
	.combout(\Mux4~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~19 .lut_mask = 16'hBBC0;
defparam \Mux4~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N25
dffeas \my_reg[14][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][27] .is_wysiwyg = "true";
defparam \my_reg[14][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N16
cycloneive_lcell_comb \Mux36~7 (
// Equation(s):
// \Mux36~7_combout  = (dcifimemload_16 & (((\my_reg[13][27]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[12][27]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[12][27]~q ),
	.datab(\my_reg[13][27]~q ),
	.datac(dcifimemload_16),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux36~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~7 .lut_mask = 16'hF0CA;
defparam \Mux36~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N24
cycloneive_lcell_comb \Mux36~8 (
// Equation(s):
// \Mux36~8_combout  = (dcifimemload_17 & ((\Mux36~7_combout  & (\my_reg[15][27]~q )) # (!\Mux36~7_combout  & ((\my_reg[14][27]~q ))))) # (!dcifimemload_17 & (((\Mux36~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[15][27]~q ),
	.datac(\my_reg[14][27]~q ),
	.datad(\Mux36~7_combout ),
	.cin(gnd),
	.combout(\Mux36~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~8 .lut_mask = 16'hDDA0;
defparam \Mux36~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N4
cycloneive_lcell_comb \my_reg[5][27]~feeder (
// Equation(s):
// \my_reg[5][27]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat6),
	.cin(gnd),
	.combout(\my_reg[5][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[5][27]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[5][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N5
dffeas \my_reg[5][27] (
	.clk(CLK),
	.d(\my_reg[5][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][27] .is_wysiwyg = "true";
defparam \my_reg[5][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N18
cycloneive_lcell_comb \Mux36~0 (
// Equation(s):
// \Mux36~0_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][27]~q ))) # (!dcifimemload_16 & (\my_reg[4][27]~q ))))

	.dataa(\my_reg[4][27]~q ),
	.datab(\my_reg[5][27]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux36~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~0 .lut_mask = 16'hFC0A;
defparam \Mux36~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N20
cycloneive_lcell_comb \Mux36~1 (
// Equation(s):
// \Mux36~1_combout  = (dcifimemload_17 & ((\Mux36~0_combout  & (\my_reg[7][27]~q )) # (!\Mux36~0_combout  & ((\my_reg[6][27]~q ))))) # (!dcifimemload_17 & (((\Mux36~0_combout ))))

	.dataa(\my_reg[7][27]~q ),
	.datab(\my_reg[6][27]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux36~0_combout ),
	.cin(gnd),
	.combout(\Mux36~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~1 .lut_mask = 16'hAFC0;
defparam \Mux36~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N23
dffeas \my_reg[11][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][27] .is_wysiwyg = "true";
defparam \my_reg[11][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N29
dffeas \my_reg[8][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][27] .is_wysiwyg = "true";
defparam \my_reg[8][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N28
cycloneive_lcell_comb \Mux36~2 (
// Equation(s):
// \Mux36~2_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\my_reg[10][27]~q )) # (!dcifimemload_17 & ((\my_reg[8][27]~q )))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[10][27]~q ),
	.datac(\my_reg[8][27]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux36~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~2 .lut_mask = 16'hEE50;
defparam \Mux36~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N22
cycloneive_lcell_comb \Mux36~3 (
// Equation(s):
// \Mux36~3_combout  = (dcifimemload_16 & ((\Mux36~2_combout  & ((\my_reg[11][27]~q ))) # (!\Mux36~2_combout  & (\my_reg[9][27]~q )))) # (!dcifimemload_16 & (((\Mux36~2_combout ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[9][27]~q ),
	.datac(\my_reg[11][27]~q ),
	.datad(\Mux36~2_combout ),
	.cin(gnd),
	.combout(\Mux36~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~3 .lut_mask = 16'hF588;
defparam \Mux36~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y42_N11
dffeas \my_reg[3][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][27] .is_wysiwyg = "true";
defparam \my_reg[3][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N10
cycloneive_lcell_comb \Mux36~4 (
// Equation(s):
// \Mux36~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][27]~q ))) # (!dcifimemload_17 & (\my_reg[1][27]~q ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[1][27]~q ),
	.datac(\my_reg[3][27]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux36~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~4 .lut_mask = 16'hA088;
defparam \Mux36~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N20
cycloneive_lcell_comb \Mux36~5 (
// Equation(s):
// \Mux36~5_combout  = (\Mux36~4_combout ) # ((!dcifimemload_16 & (\my_reg[2][27]~q  & dcifimemload_17)))

	.dataa(dcifimemload_16),
	.datab(\my_reg[2][27]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux36~4_combout ),
	.cin(gnd),
	.combout(\Mux36~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~5 .lut_mask = 16'hFF40;
defparam \Mux36~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N10
cycloneive_lcell_comb \Mux36~6 (
// Equation(s):
// \Mux36~6_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\Mux36~3_combout )) # (!dcifimemload_19 & ((\Mux36~5_combout )))))

	.dataa(dcifimemload_18),
	.datab(\Mux36~3_combout ),
	.datac(dcifimemload_19),
	.datad(\Mux36~5_combout ),
	.cin(gnd),
	.combout(\Mux36~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~6 .lut_mask = 16'hE5E0;
defparam \Mux36~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N12
cycloneive_lcell_comb \Mux36~10 (
// Equation(s):
// \Mux36~10_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[25][27]~q ))) # (!dcifimemload_19 & (\my_reg[17][27]~q ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[17][27]~q ),
	.datac(\my_reg[25][27]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux36~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~10 .lut_mask = 16'hFA44;
defparam \Mux36~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N6
cycloneive_lcell_comb \my_reg[21][27]~feeder (
// Equation(s):
// \my_reg[21][27]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat6),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[21][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][27]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[21][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N7
dffeas \my_reg[21][27] (
	.clk(CLK),
	.d(\my_reg[21][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][27] .is_wysiwyg = "true";
defparam \my_reg[21][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N22
cycloneive_lcell_comb \Mux36~11 (
// Equation(s):
// \Mux36~11_combout  = (dcifimemload_18 & ((\Mux36~10_combout  & (\my_reg[29][27]~q )) # (!\Mux36~10_combout  & ((\my_reg[21][27]~q ))))) # (!dcifimemload_18 & (((\Mux36~10_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[29][27]~q ),
	.datac(\Mux36~10_combout ),
	.datad(\my_reg[21][27]~q ),
	.cin(gnd),
	.combout(\Mux36~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~11 .lut_mask = 16'hDAD0;
defparam \Mux36~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N25
dffeas \my_reg[23][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][27] .is_wysiwyg = "true";
defparam \my_reg[23][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N24
cycloneive_lcell_comb \Mux36~17 (
// Equation(s):
// \Mux36~17_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[27][27]~q ))) # (!dcifimemload_19 & (\my_reg[19][27]~q ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[19][27]~q ),
	.datac(\my_reg[27][27]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux36~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~17 .lut_mask = 16'hFA44;
defparam \Mux36~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N24
cycloneive_lcell_comb \Mux36~18 (
// Equation(s):
// \Mux36~18_combout  = (dcifimemload_18 & ((\Mux36~17_combout  & (\my_reg[31][27]~q )) # (!\Mux36~17_combout  & ((\my_reg[23][27]~q ))))) # (!dcifimemload_18 & (((\Mux36~17_combout ))))

	.dataa(\my_reg[31][27]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[23][27]~q ),
	.datad(\Mux36~17_combout ),
	.cin(gnd),
	.combout(\Mux36~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~18 .lut_mask = 16'hBBC0;
defparam \Mux36~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y40_N19
dffeas \my_reg[24][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][27] .is_wysiwyg = "true";
defparam \my_reg[24][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N13
dffeas \my_reg[20][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][27] .is_wysiwyg = "true";
defparam \my_reg[20][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N12
cycloneive_lcell_comb \Mux36~14 (
// Equation(s):
// \Mux36~14_combout  = (dcifimemload_18 & ((dcifimemload_19) # ((\my_reg[20][27]~q )))) # (!dcifimemload_18 & (!dcifimemload_19 & ((\my_reg[16][27]~q ))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\my_reg[20][27]~q ),
	.datad(\my_reg[16][27]~q ),
	.cin(gnd),
	.combout(\Mux36~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~14 .lut_mask = 16'hB9A8;
defparam \Mux36~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N18
cycloneive_lcell_comb \Mux36~15 (
// Equation(s):
// \Mux36~15_combout  = (dcifimemload_19 & ((\Mux36~14_combout  & (\my_reg[28][27]~q )) # (!\Mux36~14_combout  & ((\my_reg[24][27]~q ))))) # (!dcifimemload_19 & (((\Mux36~14_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[28][27]~q ),
	.datac(\my_reg[24][27]~q ),
	.datad(\Mux36~14_combout ),
	.cin(gnd),
	.combout(\Mux36~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~15 .lut_mask = 16'hDDA0;
defparam \Mux36~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y42_N9
dffeas \my_reg[30][27] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][27] .is_wysiwyg = "true";
defparam \my_reg[30][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N10
cycloneive_lcell_comb \Mux36~12 (
// Equation(s):
// \Mux36~12_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\my_reg[22][27]~q )) # (!dcifimemload_18 & ((\my_reg[18][27]~q )))))

	.dataa(\my_reg[22][27]~q ),
	.datab(\my_reg[18][27]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux36~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~12 .lut_mask = 16'hFA0C;
defparam \Mux36~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N8
cycloneive_lcell_comb \Mux36~13 (
// Equation(s):
// \Mux36~13_combout  = (dcifimemload_19 & ((\Mux36~12_combout  & ((\my_reg[30][27]~q ))) # (!\Mux36~12_combout  & (\my_reg[26][27]~q )))) # (!dcifimemload_19 & (((\Mux36~12_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[26][27]~q ),
	.datac(\my_reg[30][27]~q ),
	.datad(\Mux36~12_combout ),
	.cin(gnd),
	.combout(\Mux36~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~13 .lut_mask = 16'hF588;
defparam \Mux36~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N28
cycloneive_lcell_comb \Mux36~16 (
// Equation(s):
// \Mux36~16_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux36~13_combout ))) # (!dcifimemload_17 & (\Mux36~15_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux36~15_combout ),
	.datac(dcifimemload_17),
	.datad(\Mux36~13_combout ),
	.cin(gnd),
	.combout(\Mux36~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~16 .lut_mask = 16'hF4A4;
defparam \Mux36~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N27
dffeas \my_reg[31][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][26] .is_wysiwyg = "true";
defparam \my_reg[31][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N25
dffeas \my_reg[19][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][26] .is_wysiwyg = "true";
defparam \my_reg[19][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N24
cycloneive_lcell_comb \Mux5~7 (
// Equation(s):
// \Mux5~7_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[27][26]~q )) # (!dcifimemload_24 & ((\my_reg[19][26]~q )))))

	.dataa(\my_reg[27][26]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[19][26]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux5~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~7 .lut_mask = 16'hEE30;
defparam \Mux5~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N26
cycloneive_lcell_comb \Mux5~8 (
// Equation(s):
// \Mux5~8_combout  = (dcifimemload_23 & ((\Mux5~7_combout  & ((\my_reg[31][26]~q ))) # (!\Mux5~7_combout  & (\my_reg[23][26]~q )))) # (!dcifimemload_23 & (((\Mux5~7_combout ))))

	.dataa(\my_reg[23][26]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[31][26]~q ),
	.datad(\Mux5~7_combout ),
	.cin(gnd),
	.combout(\Mux5~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~8 .lut_mask = 16'hF388;
defparam \Mux5~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N8
cycloneive_lcell_comb \my_reg[21][26]~feeder (
// Equation(s):
// \my_reg[21][26]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat7),
	.cin(gnd),
	.combout(\my_reg[21][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][26]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[21][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N9
dffeas \my_reg[21][26] (
	.clk(CLK),
	.d(\my_reg[21][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][26] .is_wysiwyg = "true";
defparam \my_reg[21][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N13
dffeas \my_reg[17][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][26] .is_wysiwyg = "true";
defparam \my_reg[17][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N12
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[25][26]~q )) # (!dcifimemload_24 & ((\my_reg[17][26]~q )))))

	.dataa(\my_reg[25][26]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[17][26]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hEE30;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N20
cycloneive_lcell_comb \my_reg[29][26]~feeder (
// Equation(s):
// \my_reg[29][26]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat7),
	.cin(gnd),
	.combout(\my_reg[29][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[29][26]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[29][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N21
dffeas \my_reg[29][26] (
	.clk(CLK),
	.d(\my_reg[29][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][26] .is_wysiwyg = "true";
defparam \my_reg[29][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N2
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// \Mux5~1_combout  = (dcifimemload_23 & ((\Mux5~0_combout  & ((\my_reg[29][26]~q ))) # (!\Mux5~0_combout  & (\my_reg[21][26]~q )))) # (!dcifimemload_23 & (((\Mux5~0_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[21][26]~q ),
	.datac(\Mux5~0_combout ),
	.datad(\my_reg[29][26]~q ),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'hF858;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N29
dffeas \my_reg[26][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][26] .is_wysiwyg = "true";
defparam \my_reg[26][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y42_N1
dffeas \my_reg[30][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][26] .is_wysiwyg = "true";
defparam \my_reg[30][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N28
cycloneive_lcell_comb \my_reg[18][26]~feeder (
// Equation(s):
// \my_reg[18][26]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat7),
	.cin(gnd),
	.combout(\my_reg[18][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[18][26]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[18][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y42_N29
dffeas \my_reg[18][26] (
	.clk(CLK),
	.d(\my_reg[18][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][26] .is_wysiwyg = "true";
defparam \my_reg[18][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N18
cycloneive_lcell_comb \Mux5~2 (
// Equation(s):
// \Mux5~2_combout  = (dcifimemload_23 & ((\my_reg[22][26]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[18][26]~q  & !dcifimemload_24))))

	.dataa(\my_reg[22][26]~q ),
	.datab(\my_reg[18][26]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~2 .lut_mask = 16'hF0AC;
defparam \Mux5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N0
cycloneive_lcell_comb \Mux5~3 (
// Equation(s):
// \Mux5~3_combout  = (dcifimemload_24 & ((\Mux5~2_combout  & ((\my_reg[30][26]~q ))) # (!\Mux5~2_combout  & (\my_reg[26][26]~q )))) # (!dcifimemload_24 & (((\Mux5~2_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[26][26]~q ),
	.datac(\my_reg[30][26]~q ),
	.datad(\Mux5~2_combout ),
	.cin(gnd),
	.combout(\Mux5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~3 .lut_mask = 16'hF588;
defparam \Mux5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N1
dffeas \my_reg[24][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][26] .is_wysiwyg = "true";
defparam \my_reg[24][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N9
dffeas \my_reg[28][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][26] .is_wysiwyg = "true";
defparam \my_reg[28][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N8
cycloneive_lcell_comb \Mux5~5 (
// Equation(s):
// \Mux5~5_combout  = (\Mux5~4_combout  & (((\my_reg[28][26]~q ) # (!dcifimemload_24)))) # (!\Mux5~4_combout  & (\my_reg[24][26]~q  & ((dcifimemload_24))))

	.dataa(\Mux5~4_combout ),
	.datab(\my_reg[24][26]~q ),
	.datac(\my_reg[28][26]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~5 .lut_mask = 16'hE4AA;
defparam \Mux5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N0
cycloneive_lcell_comb \Mux5~6 (
// Equation(s):
// \Mux5~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux5~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\Mux5~5_combout ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux5~3_combout ),
	.datad(\Mux5~5_combout ),
	.cin(gnd),
	.combout(\Mux5~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~6 .lut_mask = 16'hB9A8;
defparam \Mux5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N26
cycloneive_lcell_comb \Mux5~9 (
// Equation(s):
// \Mux5~9_combout  = (dcifimemload_21 & ((\Mux5~6_combout  & (\Mux5~8_combout )) # (!\Mux5~6_combout  & ((\Mux5~1_combout ))))) # (!dcifimemload_21 & (((\Mux5~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux5~8_combout ),
	.datac(\Mux5~1_combout ),
	.datad(\Mux5~6_combout ),
	.cin(gnd),
	.combout(\Mux5~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~9 .lut_mask = 16'hDDA0;
defparam \Mux5~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N17
dffeas \my_reg[4][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][26] .is_wysiwyg = "true";
defparam \my_reg[4][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N2
cycloneive_lcell_comb \Mux5~10 (
// Equation(s):
// \Mux5~10_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\my_reg[5][26]~q )) # (!dcifimemload_21 & ((\my_reg[4][26]~q )))))

	.dataa(\my_reg[5][26]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[4][26]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux5~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~10 .lut_mask = 16'hEE30;
defparam \Mux5~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N20
cycloneive_lcell_comb \my_reg[6][26]~feeder (
// Equation(s):
// \my_reg[6][26]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat7),
	.cin(gnd),
	.combout(\my_reg[6][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[6][26]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[6][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y43_N21
dffeas \my_reg[6][26] (
	.clk(CLK),
	.d(\my_reg[6][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][26] .is_wysiwyg = "true";
defparam \my_reg[6][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N4
cycloneive_lcell_comb \Mux5~11 (
// Equation(s):
// \Mux5~11_combout  = (\Mux5~10_combout  & ((\my_reg[7][26]~q ) # ((!dcifimemload_22)))) # (!\Mux5~10_combout  & (((dcifimemload_22 & \my_reg[6][26]~q ))))

	.dataa(\my_reg[7][26]~q ),
	.datab(\Mux5~10_combout ),
	.datac(dcifimemload_22),
	.datad(\my_reg[6][26]~q ),
	.cin(gnd),
	.combout(\Mux5~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~11 .lut_mask = 16'hBC8C;
defparam \Mux5~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N11
dffeas \my_reg[11][26] (
	.clk(CLK),
	.d(wdat7),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][26] .is_wysiwyg = "true";
defparam \my_reg[11][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N16
cycloneive_lcell_comb \my_reg[10][26]~feeder (
// Equation(s):
// \my_reg[10][26]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat7),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[10][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[10][26]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[10][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y38_N17
dffeas \my_reg[10][26] (
	.clk(CLK),
	.d(\my_reg[10][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][26] .is_wysiwyg = "true";
defparam \my_reg[10][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N21
dffeas \my_reg[8][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][26] .is_wysiwyg = "true";
defparam \my_reg[8][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N20
cycloneive_lcell_comb \Mux5~12 (
// Equation(s):
// \Mux5~12_combout  = (dcifimemload_22 & ((\my_reg[10][26]~q ) # ((dcifimemload_21)))) # (!dcifimemload_22 & (((\my_reg[8][26]~q  & !dcifimemload_21))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[10][26]~q ),
	.datac(\my_reg[8][26]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux5~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~12 .lut_mask = 16'hAAD8;
defparam \Mux5~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N24
cycloneive_lcell_comb \Mux5~13 (
// Equation(s):
// \Mux5~13_combout  = (\Mux5~12_combout  & (((\my_reg[11][26]~q ) # (!dcifimemload_21)))) # (!\Mux5~12_combout  & (\my_reg[9][26]~q  & ((dcifimemload_21))))

	.dataa(\my_reg[9][26]~q ),
	.datab(\my_reg[11][26]~q ),
	.datac(\Mux5~12_combout ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux5~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~13 .lut_mask = 16'hCAF0;
defparam \Mux5~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y42_N23
dffeas \my_reg[3][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][26] .is_wysiwyg = "true";
defparam \my_reg[3][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y42_N1
dffeas \my_reg[1][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][26] .is_wysiwyg = "true";
defparam \my_reg[1][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N0
cycloneive_lcell_comb \Mux5~14 (
// Equation(s):
// \Mux5~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\my_reg[3][26]~q )) # (!dcifimemload_22 & ((\my_reg[1][26]~q )))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[3][26]~q ),
	.datac(\my_reg[1][26]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux5~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~14 .lut_mask = 16'h88A0;
defparam \Mux5~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N30
cycloneive_lcell_comb \Mux5~15 (
// Equation(s):
// \Mux5~15_combout  = (\Mux5~14_combout ) # ((\my_reg[2][26]~q  & (!dcifimemload_21 & dcifimemload_22)))

	.dataa(\my_reg[2][26]~q ),
	.datab(dcifimemload_21),
	.datac(dcifimemload_22),
	.datad(\Mux5~14_combout ),
	.cin(gnd),
	.combout(\Mux5~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~15 .lut_mask = 16'hFF20;
defparam \Mux5~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N8
cycloneive_lcell_comb \Mux5~16 (
// Equation(s):
// \Mux5~16_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\Mux5~13_combout )) # (!dcifimemload_24 & ((\Mux5~15_combout )))))

	.dataa(dcifimemload_23),
	.datab(\Mux5~13_combout ),
	.datac(\Mux5~15_combout ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux5~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~16 .lut_mask = 16'hEE50;
defparam \Mux5~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N26
cycloneive_lcell_comb \my_reg[15][26]~feeder (
// Equation(s):
// \my_reg[15][26]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat7),
	.cin(gnd),
	.combout(\my_reg[15][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[15][26]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[15][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N27
dffeas \my_reg[15][26] (
	.clk(CLK),
	.d(\my_reg[15][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][26] .is_wysiwyg = "true";
defparam \my_reg[15][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N19
dffeas \my_reg[13][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][26] .is_wysiwyg = "true";
defparam \my_reg[13][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N31
dffeas \my_reg[12][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][26] .is_wysiwyg = "true";
defparam \my_reg[12][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N30
cycloneive_lcell_comb \Mux5~17 (
// Equation(s):
// \Mux5~17_combout  = (dcifimemload_21 & ((\my_reg[13][26]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][26]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[13][26]~q ),
	.datac(\my_reg[12][26]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux5~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~17 .lut_mask = 16'hAAD8;
defparam \Mux5~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N10
cycloneive_lcell_comb \Mux5~18 (
// Equation(s):
// \Mux5~18_combout  = (\Mux5~17_combout  & (((\my_reg[15][26]~q ) # (!dcifimemload_22)))) # (!\Mux5~17_combout  & (\my_reg[14][26]~q  & ((dcifimemload_22))))

	.dataa(\my_reg[14][26]~q ),
	.datab(\my_reg[15][26]~q ),
	.datac(\Mux5~17_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux5~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~18 .lut_mask = 16'hCAF0;
defparam \Mux5~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N16
cycloneive_lcell_comb \Mux5~19 (
// Equation(s):
// \Mux5~19_combout  = (dcifimemload_23 & ((\Mux5~16_combout  & ((\Mux5~18_combout ))) # (!\Mux5~16_combout  & (\Mux5~11_combout )))) # (!dcifimemload_23 & (((\Mux5~16_combout ))))

	.dataa(dcifimemload_23),
	.datab(\Mux5~11_combout ),
	.datac(\Mux5~16_combout ),
	.datad(\Mux5~18_combout ),
	.cin(gnd),
	.combout(\Mux5~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~19 .lut_mask = 16'hF858;
defparam \Mux5~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N5
dffeas \my_reg[14][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][26] .is_wysiwyg = "true";
defparam \my_reg[14][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N18
cycloneive_lcell_comb \Mux37~7 (
// Equation(s):
// \Mux37~7_combout  = (dcifimemload_16 & (((\my_reg[13][26]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[12][26]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[12][26]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[13][26]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux37~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~7 .lut_mask = 16'hCCE2;
defparam \Mux37~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N4
cycloneive_lcell_comb \Mux37~8 (
// Equation(s):
// \Mux37~8_combout  = (dcifimemload_17 & ((\Mux37~7_combout  & (\my_reg[15][26]~q )) # (!\Mux37~7_combout  & ((\my_reg[14][26]~q ))))) # (!dcifimemload_17 & (((\Mux37~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[15][26]~q ),
	.datac(\my_reg[14][26]~q ),
	.datad(\Mux37~7_combout ),
	.cin(gnd),
	.combout(\Mux37~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~8 .lut_mask = 16'hDDA0;
defparam \Mux37~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N6
cycloneive_lcell_comb \my_reg[9][26]~feeder (
// Equation(s):
// \my_reg[9][26]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat7),
	.cin(gnd),
	.combout(\my_reg[9][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[9][26]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[9][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y43_N7
dffeas \my_reg[9][26] (
	.clk(CLK),
	.d(\my_reg[9][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][26] .is_wysiwyg = "true";
defparam \my_reg[9][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N18
cycloneive_lcell_comb \Mux37~0 (
// Equation(s):
// \Mux37~0_combout  = (dcifimemload_17 & (((\my_reg[10][26]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\my_reg[8][26]~q  & ((!dcifimemload_16))))

	.dataa(\my_reg[8][26]~q ),
	.datab(\my_reg[10][26]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~0 .lut_mask = 16'hF0CA;
defparam \Mux37~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N4
cycloneive_lcell_comb \Mux37~1 (
// Equation(s):
// \Mux37~1_combout  = (dcifimemload_16 & ((\Mux37~0_combout  & (\my_reg[11][26]~q )) # (!\Mux37~0_combout  & ((\my_reg[9][26]~q ))))) # (!dcifimemload_16 & (((\Mux37~0_combout ))))

	.dataa(\my_reg[11][26]~q ),
	.datab(\my_reg[9][26]~q ),
	.datac(dcifimemload_16),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\Mux37~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~1 .lut_mask = 16'hAFC0;
defparam \Mux37~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N22
cycloneive_lcell_comb \Mux37~4 (
// Equation(s):
// \Mux37~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][26]~q ))) # (!dcifimemload_17 & (\my_reg[1][26]~q ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[1][26]~q ),
	.datac(\my_reg[3][26]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux37~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~4 .lut_mask = 16'hA088;
defparam \Mux37~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N8
cycloneive_lcell_comb \Mux37~5 (
// Equation(s):
// \Mux37~5_combout  = (\Mux37~4_combout ) # ((\my_reg[2][26]~q  & (dcifimemload_17 & !dcifimemload_16)))

	.dataa(\my_reg[2][26]~q ),
	.datab(dcifimemload_17),
	.datac(\Mux37~4_combout ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux37~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~5 .lut_mask = 16'hF0F8;
defparam \Mux37~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N19
dffeas \my_reg[7][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][26] .is_wysiwyg = "true";
defparam \my_reg[7][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N4
cycloneive_lcell_comb \my_reg[5][26]~feeder (
// Equation(s):
// \my_reg[5][26]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat7),
	.cin(gnd),
	.combout(\my_reg[5][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[5][26]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[5][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y43_N5
dffeas \my_reg[5][26] (
	.clk(CLK),
	.d(\my_reg[5][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][26] .is_wysiwyg = "true";
defparam \my_reg[5][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N16
cycloneive_lcell_comb \Mux37~2 (
// Equation(s):
// \Mux37~2_combout  = (dcifimemload_16 & ((\my_reg[5][26]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\my_reg[4][26]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[5][26]~q ),
	.datac(\my_reg[4][26]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux37~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~2 .lut_mask = 16'hAAD8;
defparam \Mux37~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N18
cycloneive_lcell_comb \Mux37~3 (
// Equation(s):
// \Mux37~3_combout  = (dcifimemload_17 & ((\Mux37~2_combout  & ((\my_reg[7][26]~q ))) # (!\Mux37~2_combout  & (\my_reg[6][26]~q )))) # (!dcifimemload_17 & (((\Mux37~2_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[6][26]~q ),
	.datac(\my_reg[7][26]~q ),
	.datad(\Mux37~2_combout ),
	.cin(gnd),
	.combout(\Mux37~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~3 .lut_mask = 16'hF588;
defparam \Mux37~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N26
cycloneive_lcell_comb \Mux37~6 (
// Equation(s):
// \Mux37~6_combout  = (dcifimemload_18 & ((dcifimemload_19) # ((\Mux37~3_combout )))) # (!dcifimemload_18 & (!dcifimemload_19 & (\Mux37~5_combout )))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux37~5_combout ),
	.datad(\Mux37~3_combout ),
	.cin(gnd),
	.combout(\Mux37~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~6 .lut_mask = 16'hBA98;
defparam \Mux37~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N0
cycloneive_lcell_comb \my_reg[27][26]~feeder (
// Equation(s):
// \my_reg[27][26]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat7),
	.cin(gnd),
	.combout(\my_reg[27][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[27][26]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[27][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N1
dffeas \my_reg[27][26] (
	.clk(CLK),
	.d(\my_reg[27][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][26] .is_wysiwyg = "true";
defparam \my_reg[27][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N0
cycloneive_lcell_comb \Mux37~17 (
// Equation(s):
// \Mux37~17_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\my_reg[23][26]~q )) # (!dcifimemload_18 & ((\my_reg[19][26]~q )))))

	.dataa(\my_reg[23][26]~q ),
	.datab(\my_reg[19][26]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux37~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~17 .lut_mask = 16'hFA0C;
defparam \Mux37~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N18
cycloneive_lcell_comb \Mux37~18 (
// Equation(s):
// \Mux37~18_combout  = (dcifimemload_19 & ((\Mux37~17_combout  & (\my_reg[31][26]~q )) # (!\Mux37~17_combout  & ((\my_reg[27][26]~q ))))) # (!dcifimemload_19 & (((\Mux37~17_combout ))))

	.dataa(\my_reg[31][26]~q ),
	.datab(\my_reg[27][26]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux37~17_combout ),
	.cin(gnd),
	.combout(\Mux37~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~18 .lut_mask = 16'hAFC0;
defparam \Mux37~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N30
cycloneive_lcell_comb \my_reg[25][26]~feeder (
// Equation(s):
// \my_reg[25][26]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat7),
	.cin(gnd),
	.combout(\my_reg[25][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][26]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[25][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N31
dffeas \my_reg[25][26] (
	.clk(CLK),
	.d(\my_reg[25][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][26] .is_wysiwyg = "true";
defparam \my_reg[25][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N28
cycloneive_lcell_comb \Mux37~10 (
// Equation(s):
// \Mux37~10_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[21][26]~q ))) # (!dcifimemload_18 & (\my_reg[17][26]~q ))))

	.dataa(\my_reg[17][26]~q ),
	.datab(\my_reg[21][26]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux37~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~10 .lut_mask = 16'hFC0A;
defparam \Mux37~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N14
cycloneive_lcell_comb \Mux37~11 (
// Equation(s):
// \Mux37~11_combout  = (dcifimemload_19 & ((\Mux37~10_combout  & ((\my_reg[29][26]~q ))) # (!\Mux37~10_combout  & (\my_reg[25][26]~q )))) # (!dcifimemload_19 & (((\Mux37~10_combout ))))

	.dataa(\my_reg[25][26]~q ),
	.datab(\my_reg[29][26]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux37~10_combout ),
	.cin(gnd),
	.combout(\Mux37~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~11 .lut_mask = 16'hCFA0;
defparam \Mux37~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N3
dffeas \my_reg[20][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][26] .is_wysiwyg = "true";
defparam \my_reg[20][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N31
dffeas \my_reg[16][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][26] .is_wysiwyg = "true";
defparam \my_reg[16][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N0
cycloneive_lcell_comb \Mux37~14 (
// Equation(s):
// \Mux37~14_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & (\my_reg[24][26]~q )) # (!dcifimemload_19 & ((\my_reg[16][26]~q )))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\my_reg[24][26]~q ),
	.datad(\my_reg[16][26]~q ),
	.cin(gnd),
	.combout(\Mux37~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~14 .lut_mask = 16'hD9C8;
defparam \Mux37~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N2
cycloneive_lcell_comb \Mux37~15 (
// Equation(s):
// \Mux37~15_combout  = (dcifimemload_18 & ((\Mux37~14_combout  & (\my_reg[28][26]~q )) # (!\Mux37~14_combout  & ((\my_reg[20][26]~q ))))) # (!dcifimemload_18 & (((\Mux37~14_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[28][26]~q ),
	.datac(\my_reg[20][26]~q ),
	.datad(\Mux37~14_combout ),
	.cin(gnd),
	.combout(\Mux37~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~15 .lut_mask = 16'hDDA0;
defparam \Mux37~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N7
dffeas \my_reg[22][26] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][26] .is_wysiwyg = "true";
defparam \my_reg[22][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N28
cycloneive_lcell_comb \Mux37~12 (
// Equation(s):
// \Mux37~12_combout  = (dcifimemload_19 & (((\my_reg[26][26]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[18][26]~q  & ((!dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[18][26]~q ),
	.datac(\my_reg[26][26]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux37~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~12 .lut_mask = 16'hAAE4;
defparam \Mux37~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N6
cycloneive_lcell_comb \Mux37~13 (
// Equation(s):
// \Mux37~13_combout  = (dcifimemload_18 & ((\Mux37~12_combout  & (\my_reg[30][26]~q )) # (!\Mux37~12_combout  & ((\my_reg[22][26]~q ))))) # (!dcifimemload_18 & (((\Mux37~12_combout ))))

	.dataa(\my_reg[30][26]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[22][26]~q ),
	.datad(\Mux37~12_combout ),
	.cin(gnd),
	.combout(\Mux37~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~13 .lut_mask = 16'hBBC0;
defparam \Mux37~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N6
cycloneive_lcell_comb \Mux37~16 (
// Equation(s):
// \Mux37~16_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux37~13_combout ))) # (!dcifimemload_17 & (\Mux37~15_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux37~15_combout ),
	.datac(dcifimemload_17),
	.datad(\Mux37~13_combout ),
	.cin(gnd),
	.combout(\Mux37~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~16 .lut_mask = 16'hF4A4;
defparam \Mux37~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y42_N19
dffeas \my_reg[9][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][25] .is_wysiwyg = "true";
defparam \my_reg[9][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N15
dffeas \my_reg[11][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][25] .is_wysiwyg = "true";
defparam \my_reg[11][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y42_N21
dffeas \my_reg[10][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][25] .is_wysiwyg = "true";
defparam \my_reg[10][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N29
dffeas \my_reg[8][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][25] .is_wysiwyg = "true";
defparam \my_reg[8][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N28
cycloneive_lcell_comb \Mux6~10 (
// Equation(s):
// \Mux6~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][25]~q )) # (!dcifimemload_22 & ((\my_reg[8][25]~q )))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[10][25]~q ),
	.datac(\my_reg[8][25]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux6~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~10 .lut_mask = 16'hEE50;
defparam \Mux6~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N14
cycloneive_lcell_comb \Mux6~11 (
// Equation(s):
// \Mux6~11_combout  = (dcifimemload_21 & ((\Mux6~10_combout  & ((\my_reg[11][25]~q ))) # (!\Mux6~10_combout  & (\my_reg[9][25]~q )))) # (!dcifimemload_21 & (((\Mux6~10_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][25]~q ),
	.datac(\my_reg[11][25]~q ),
	.datad(\Mux6~10_combout ),
	.cin(gnd),
	.combout(\Mux6~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~11 .lut_mask = 16'hF588;
defparam \Mux6~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N5
dffeas \my_reg[14][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][25] .is_wysiwyg = "true";
defparam \my_reg[14][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N7
dffeas \my_reg[15][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][25] .is_wysiwyg = "true";
defparam \my_reg[15][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N13
dffeas \my_reg[13][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][25] .is_wysiwyg = "true";
defparam \my_reg[13][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N13
dffeas \my_reg[12][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][25] .is_wysiwyg = "true";
defparam \my_reg[12][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N12
cycloneive_lcell_comb \Mux6~17 (
// Equation(s):
// \Mux6~17_combout  = (dcifimemload_21 & ((\my_reg[13][25]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][25]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[13][25]~q ),
	.datac(\my_reg[12][25]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux6~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~17 .lut_mask = 16'hAAD8;
defparam \Mux6~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N6
cycloneive_lcell_comb \Mux6~18 (
// Equation(s):
// \Mux6~18_combout  = (dcifimemload_22 & ((\Mux6~17_combout  & ((\my_reg[15][25]~q ))) # (!\Mux6~17_combout  & (\my_reg[14][25]~q )))) # (!dcifimemload_22 & (((\Mux6~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[14][25]~q ),
	.datac(\my_reg[15][25]~q ),
	.datad(\Mux6~17_combout ),
	.cin(gnd),
	.combout(\Mux6~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~18 .lut_mask = 16'hF588;
defparam \Mux6~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N1
dffeas \my_reg[6][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][25] .is_wysiwyg = "true";
defparam \my_reg[6][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y43_N7
dffeas \my_reg[7][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][25] .is_wysiwyg = "true";
defparam \my_reg[7][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y43_N1
dffeas \my_reg[4][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][25] .is_wysiwyg = "true";
defparam \my_reg[4][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y42_N23
dffeas \my_reg[5][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][25] .is_wysiwyg = "true";
defparam \my_reg[5][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N0
cycloneive_lcell_comb \Mux6~12 (
// Equation(s):
// \Mux6~12_combout  = (dcifimemload_22 & (dcifimemload_21)) # (!dcifimemload_22 & ((dcifimemload_21 & ((\my_reg[5][25]~q ))) # (!dcifimemload_21 & (\my_reg[4][25]~q ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\my_reg[4][25]~q ),
	.datad(\my_reg[5][25]~q ),
	.cin(gnd),
	.combout(\Mux6~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~12 .lut_mask = 16'hDC98;
defparam \Mux6~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N6
cycloneive_lcell_comb \Mux6~13 (
// Equation(s):
// \Mux6~13_combout  = (dcifimemload_22 & ((\Mux6~12_combout  & ((\my_reg[7][25]~q ))) # (!\Mux6~12_combout  & (\my_reg[6][25]~q )))) # (!dcifimemload_22 & (((\Mux6~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[6][25]~q ),
	.datac(\my_reg[7][25]~q ),
	.datad(\Mux6~12_combout ),
	.cin(gnd),
	.combout(\Mux6~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~13 .lut_mask = 16'hF588;
defparam \Mux6~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N11
dffeas \my_reg[2][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][25] .is_wysiwyg = "true";
defparam \my_reg[2][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N10
cycloneive_lcell_comb \Mux6~15 (
// Equation(s):
// \Mux6~15_combout  = (\Mux6~14_combout ) # ((dcifimemload_22 & (\my_reg[2][25]~q  & !dcifimemload_21)))

	.dataa(\Mux6~14_combout ),
	.datab(dcifimemload_22),
	.datac(\my_reg[2][25]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux6~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~15 .lut_mask = 16'hAAEA;
defparam \Mux6~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N20
cycloneive_lcell_comb \Mux6~16 (
// Equation(s):
// \Mux6~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & (\Mux6~13_combout )) # (!dcifimemload_23 & ((\Mux6~15_combout )))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux6~13_combout ),
	.datad(\Mux6~15_combout ),
	.cin(gnd),
	.combout(\Mux6~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~16 .lut_mask = 16'hD9C8;
defparam \Mux6~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N14
cycloneive_lcell_comb \Mux6~19 (
// Equation(s):
// \Mux6~19_combout  = (dcifimemload_24 & ((\Mux6~16_combout  & ((\Mux6~18_combout ))) # (!\Mux6~16_combout  & (\Mux6~11_combout )))) # (!dcifimemload_24 & (((\Mux6~16_combout ))))

	.dataa(dcifimemload_24),
	.datab(\Mux6~11_combout ),
	.datac(\Mux6~18_combout ),
	.datad(\Mux6~16_combout ),
	.cin(gnd),
	.combout(\Mux6~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~19 .lut_mask = 16'hF588;
defparam \Mux6~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N5
dffeas \my_reg[29][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][25] .is_wysiwyg = "true";
defparam \my_reg[29][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N5
dffeas \my_reg[25][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][25] .is_wysiwyg = "true";
defparam \my_reg[25][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N3
dffeas \my_reg[17][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][25] .is_wysiwyg = "true";
defparam \my_reg[17][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N2
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (dcifimemload_23 & ((\my_reg[21][25]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[17][25]~q  & !dcifimemload_24))))

	.dataa(\my_reg[21][25]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[17][25]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'hCCB8;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N4
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// \Mux6~1_combout  = (dcifimemload_24 & ((\Mux6~0_combout  & (\my_reg[29][25]~q )) # (!\Mux6~0_combout  & ((\my_reg[25][25]~q ))))) # (!dcifimemload_24 & (((\Mux6~0_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[29][25]~q ),
	.datac(\my_reg[25][25]~q ),
	.datad(\Mux6~0_combout ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hDDA0;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y42_N17
dffeas \my_reg[20][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][25] .is_wysiwyg = "true";
defparam \my_reg[20][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N17
dffeas \my_reg[28][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][25] .is_wysiwyg = "true";
defparam \my_reg[28][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y42_N31
dffeas \my_reg[24][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][25] .is_wysiwyg = "true";
defparam \my_reg[24][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N3
dffeas \my_reg[16][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][25] .is_wysiwyg = "true";
defparam \my_reg[16][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N2
cycloneive_lcell_comb \Mux6~4 (
// Equation(s):
// \Mux6~4_combout  = (dcifimemload_24 & ((\my_reg[24][25]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\my_reg[16][25]~q  & !dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[24][25]~q ),
	.datac(\my_reg[16][25]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux6~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~4 .lut_mask = 16'hAAD8;
defparam \Mux6~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N16
cycloneive_lcell_comb \Mux6~5 (
// Equation(s):
// \Mux6~5_combout  = (dcifimemload_23 & ((\Mux6~4_combout  & ((\my_reg[28][25]~q ))) # (!\Mux6~4_combout  & (\my_reg[20][25]~q )))) # (!dcifimemload_23 & (((\Mux6~4_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[20][25]~q ),
	.datac(\my_reg[28][25]~q ),
	.datad(\Mux6~4_combout ),
	.cin(gnd),
	.combout(\Mux6~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~5 .lut_mask = 16'hF588;
defparam \Mux6~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y42_N31
dffeas \my_reg[30][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][25] .is_wysiwyg = "true";
defparam \my_reg[30][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y42_N27
dffeas \my_reg[26][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][25] .is_wysiwyg = "true";
defparam \my_reg[26][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N24
cycloneive_lcell_comb \Mux6~2 (
// Equation(s):
// \Mux6~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\my_reg[26][25]~q ))) # (!dcifimemload_24 & (\my_reg[18][25]~q ))))

	.dataa(\my_reg[18][25]~q ),
	.datab(\my_reg[26][25]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~2 .lut_mask = 16'hFC0A;
defparam \Mux6~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N30
cycloneive_lcell_comb \Mux6~3 (
// Equation(s):
// \Mux6~3_combout  = (dcifimemload_23 & ((\Mux6~2_combout  & ((\my_reg[30][25]~q ))) # (!\Mux6~2_combout  & (\my_reg[22][25]~q )))) # (!dcifimemload_23 & (((\Mux6~2_combout ))))

	.dataa(\my_reg[22][25]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[30][25]~q ),
	.datad(\Mux6~2_combout ),
	.cin(gnd),
	.combout(\Mux6~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~3 .lut_mask = 16'hF388;
defparam \Mux6~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N8
cycloneive_lcell_comb \Mux6~6 (
// Equation(s):
// \Mux6~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux6~3_combout ))) # (!dcifimemload_22 & (\Mux6~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux6~5_combout ),
	.datad(\Mux6~3_combout ),
	.cin(gnd),
	.combout(\Mux6~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~6 .lut_mask = 16'hDC98;
defparam \Mux6~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N3
dffeas \my_reg[27][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][25] .is_wysiwyg = "true";
defparam \my_reg[27][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N7
dffeas \my_reg[31][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][25] .is_wysiwyg = "true";
defparam \my_reg[31][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N21
dffeas \my_reg[23][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][25] .is_wysiwyg = "true";
defparam \my_reg[23][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N20
cycloneive_lcell_comb \Mux6~7 (
// Equation(s):
// \Mux6~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\my_reg[23][25]~q ))) # (!dcifimemload_23 & (\my_reg[19][25]~q ))))

	.dataa(\my_reg[19][25]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[23][25]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux6~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~7 .lut_mask = 16'hFC22;
defparam \Mux6~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N6
cycloneive_lcell_comb \Mux6~8 (
// Equation(s):
// \Mux6~8_combout  = (dcifimemload_24 & ((\Mux6~7_combout  & ((\my_reg[31][25]~q ))) # (!\Mux6~7_combout  & (\my_reg[27][25]~q )))) # (!dcifimemload_24 & (((\Mux6~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[27][25]~q ),
	.datac(\my_reg[31][25]~q ),
	.datad(\Mux6~7_combout ),
	.cin(gnd),
	.combout(\Mux6~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~8 .lut_mask = 16'hF588;
defparam \Mux6~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N6
cycloneive_lcell_comb \Mux6~9 (
// Equation(s):
// \Mux6~9_combout  = (dcifimemload_21 & ((\Mux6~6_combout  & ((\Mux6~8_combout ))) # (!\Mux6~6_combout  & (\Mux6~1_combout )))) # (!dcifimemload_21 & (((\Mux6~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux6~1_combout ),
	.datac(\Mux6~6_combout ),
	.datad(\Mux6~8_combout ),
	.cin(gnd),
	.combout(\Mux6~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~9 .lut_mask = 16'hF858;
defparam \Mux6~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N29
dffeas \my_reg[3][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][25] .is_wysiwyg = "true";
defparam \my_reg[3][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N28
cycloneive_lcell_comb \Mux38~4 (
// Equation(s):
// \Mux38~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][25]~q ))) # (!dcifimemload_17 & (\my_reg[1][25]~q ))))

	.dataa(\my_reg[1][25]~q ),
	.datab(dcifimemload_17),
	.datac(\my_reg[3][25]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux38~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~4 .lut_mask = 16'hE200;
defparam \Mux38~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N8
cycloneive_lcell_comb \Mux38~5 (
// Equation(s):
// \Mux38~5_combout  = (\Mux38~4_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \my_reg[2][25]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\my_reg[2][25]~q ),
	.datad(\Mux38~4_combout ),
	.cin(gnd),
	.combout(\Mux38~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~5 .lut_mask = 16'hFF20;
defparam \Mux38~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N20
cycloneive_lcell_comb \Mux38~2 (
// Equation(s):
// \Mux38~2_combout  = (dcifimemload_17 & (((\my_reg[10][25]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\my_reg[8][25]~q  & ((!dcifimemload_16))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[8][25]~q ),
	.datac(\my_reg[10][25]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux38~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~2 .lut_mask = 16'hAAE4;
defparam \Mux38~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N18
cycloneive_lcell_comb \Mux38~3 (
// Equation(s):
// \Mux38~3_combout  = (\Mux38~2_combout  & ((\my_reg[11][25]~q ) # ((!dcifimemload_16)))) # (!\Mux38~2_combout  & (((\my_reg[9][25]~q  & dcifimemload_16))))

	.dataa(\my_reg[11][25]~q ),
	.datab(\Mux38~2_combout ),
	.datac(\my_reg[9][25]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux38~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~3 .lut_mask = 16'hB8CC;
defparam \Mux38~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N26
cycloneive_lcell_comb \Mux38~6 (
// Equation(s):
// \Mux38~6_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\Mux38~3_combout )))) # (!dcifimemload_19 & (!dcifimemload_18 & (\Mux38~5_combout )))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux38~5_combout ),
	.datad(\Mux38~3_combout ),
	.cin(gnd),
	.combout(\Mux38~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~6 .lut_mask = 16'hBA98;
defparam \Mux38~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N12
cycloneive_lcell_comb \Mux38~7 (
// Equation(s):
// \Mux38~7_combout  = (dcifimemload_16 & (((\my_reg[13][25]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[12][25]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[12][25]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[13][25]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux38~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~7 .lut_mask = 16'hCCE2;
defparam \Mux38~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N4
cycloneive_lcell_comb \Mux38~8 (
// Equation(s):
// \Mux38~8_combout  = (dcifimemload_17 & ((\Mux38~7_combout  & (\my_reg[15][25]~q )) # (!\Mux38~7_combout  & ((\my_reg[14][25]~q ))))) # (!dcifimemload_17 & (((\Mux38~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[15][25]~q ),
	.datac(\my_reg[14][25]~q ),
	.datad(\Mux38~7_combout ),
	.cin(gnd),
	.combout(\Mux38~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~8 .lut_mask = 16'hDDA0;
defparam \Mux38~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N22
cycloneive_lcell_comb \Mux38~0 (
// Equation(s):
// \Mux38~0_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][25]~q ))) # (!dcifimemload_16 & (\my_reg[4][25]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[4][25]~q ),
	.datac(\my_reg[5][25]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux38~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~0 .lut_mask = 16'hFA44;
defparam \Mux38~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N0
cycloneive_lcell_comb \Mux38~1 (
// Equation(s):
// \Mux38~1_combout  = (\Mux38~0_combout  & ((\my_reg[7][25]~q ) # ((!dcifimemload_17)))) # (!\Mux38~0_combout  & (((\my_reg[6][25]~q  & dcifimemload_17))))

	.dataa(\Mux38~0_combout ),
	.datab(\my_reg[7][25]~q ),
	.datac(\my_reg[6][25]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux38~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~1 .lut_mask = 16'hD8AA;
defparam \Mux38~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N30
cycloneive_lcell_comb \my_reg[21][25]~feeder (
// Equation(s):
// \my_reg[21][25]~feeder_combout  = \wdat~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat8),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[21][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][25]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[21][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N31
dffeas \my_reg[21][25] (
	.clk(CLK),
	.d(\my_reg[21][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][25] .is_wysiwyg = "true";
defparam \my_reg[21][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N4
cycloneive_lcell_comb \Mux38~10 (
// Equation(s):
// \Mux38~10_combout  = (dcifimemload_19 & (((\my_reg[25][25]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[17][25]~q  & ((!dcifimemload_18))))

	.dataa(\my_reg[17][25]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[25][25]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux38~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~10 .lut_mask = 16'hCCE2;
defparam \Mux38~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N4
cycloneive_lcell_comb \Mux38~11 (
// Equation(s):
// \Mux38~11_combout  = (\Mux38~10_combout  & (((\my_reg[29][25]~q ) # (!dcifimemload_18)))) # (!\Mux38~10_combout  & (\my_reg[21][25]~q  & ((dcifimemload_18))))

	.dataa(\my_reg[21][25]~q ),
	.datab(\Mux38~10_combout ),
	.datac(\my_reg[29][25]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux38~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~11 .lut_mask = 16'hE2CC;
defparam \Mux38~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N24
cycloneive_lcell_comb \my_reg[19][25]~feeder (
// Equation(s):
// \my_reg[19][25]~feeder_combout  = \wdat~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat8),
	.cin(gnd),
	.combout(\my_reg[19][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[19][25]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[19][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y33_N25
dffeas \my_reg[19][25] (
	.clk(CLK),
	.d(\my_reg[19][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][25] .is_wysiwyg = "true";
defparam \my_reg[19][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N2
cycloneive_lcell_comb \Mux38~17 (
// Equation(s):
// \Mux38~17_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[27][25]~q ))) # (!dcifimemload_19 & (\my_reg[19][25]~q ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[19][25]~q ),
	.datac(\my_reg[27][25]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux38~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~17 .lut_mask = 16'hFA44;
defparam \Mux38~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N16
cycloneive_lcell_comb \Mux38~18 (
// Equation(s):
// \Mux38~18_combout  = (\Mux38~17_combout  & ((\my_reg[31][25]~q ) # ((!dcifimemload_18)))) # (!\Mux38~17_combout  & (((\my_reg[23][25]~q  & dcifimemload_18))))

	.dataa(\my_reg[31][25]~q ),
	.datab(\my_reg[23][25]~q ),
	.datac(\Mux38~17_combout ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux38~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~18 .lut_mask = 16'hACF0;
defparam \Mux38~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N16
cycloneive_lcell_comb \Mux38~14 (
// Equation(s):
// \Mux38~14_combout  = (dcifimemload_18 & (((\my_reg[20][25]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[16][25]~q  & ((!dcifimemload_19))))

	.dataa(\my_reg[16][25]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[20][25]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux38~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~14 .lut_mask = 16'hCCE2;
defparam \Mux38~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N30
cycloneive_lcell_comb \Mux38~15 (
// Equation(s):
// \Mux38~15_combout  = (dcifimemload_19 & ((\Mux38~14_combout  & (\my_reg[28][25]~q )) # (!\Mux38~14_combout  & ((\my_reg[24][25]~q ))))) # (!dcifimemload_19 & (((\Mux38~14_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[28][25]~q ),
	.datac(\my_reg[24][25]~q ),
	.datad(\Mux38~14_combout ),
	.cin(gnd),
	.combout(\Mux38~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~15 .lut_mask = 16'hDDA0;
defparam \Mux38~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N6
cycloneive_lcell_comb \my_reg[18][25]~feeder (
// Equation(s):
// \my_reg[18][25]~feeder_combout  = \wdat~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat8),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[18][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[18][25]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[18][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y42_N7
dffeas \my_reg[18][25] (
	.clk(CLK),
	.d(\my_reg[18][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][25] .is_wysiwyg = "true";
defparam \my_reg[18][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y42_N5
dffeas \my_reg[22][25] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][25] .is_wysiwyg = "true";
defparam \my_reg[22][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N4
cycloneive_lcell_comb \Mux38~12 (
// Equation(s):
// \Mux38~12_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[22][25]~q ))) # (!dcifimemload_18 & (\my_reg[18][25]~q ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[18][25]~q ),
	.datac(\my_reg[22][25]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux38~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~12 .lut_mask = 16'hFA44;
defparam \Mux38~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N26
cycloneive_lcell_comb \Mux38~13 (
// Equation(s):
// \Mux38~13_combout  = (dcifimemload_19 & ((\Mux38~12_combout  & (\my_reg[30][25]~q )) # (!\Mux38~12_combout  & ((\my_reg[26][25]~q ))))) # (!dcifimemload_19 & (((\Mux38~12_combout ))))

	.dataa(\my_reg[30][25]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[26][25]~q ),
	.datad(\Mux38~12_combout ),
	.cin(gnd),
	.combout(\Mux38~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~13 .lut_mask = 16'hBBC0;
defparam \Mux38~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N12
cycloneive_lcell_comb \Mux38~16 (
// Equation(s):
// \Mux38~16_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux38~13_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & (\Mux38~15_combout )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux38~15_combout ),
	.datad(\Mux38~13_combout ),
	.cin(gnd),
	.combout(\Mux38~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~16 .lut_mask = 16'hBA98;
defparam \Mux38~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N4
cycloneive_lcell_comb \my_reg[21][24]~feeder (
// Equation(s):
// \my_reg[21][24]~feeder_combout  = \wdat~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat9),
	.cin(gnd),
	.combout(\my_reg[21][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][24]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[21][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N5
dffeas \my_reg[21][24] (
	.clk(CLK),
	.d(\my_reg[21][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][24] .is_wysiwyg = "true";
defparam \my_reg[21][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N31
dffeas \my_reg[29][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][24] .is_wysiwyg = "true";
defparam \my_reg[29][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N8
cycloneive_lcell_comb \my_reg[25][24]~feeder (
// Equation(s):
// \my_reg[25][24]~feeder_combout  = \wdat~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat9),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[25][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][24]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[25][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N9
dffeas \my_reg[25][24] (
	.clk(CLK),
	.d(\my_reg[25][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][24] .is_wysiwyg = "true";
defparam \my_reg[25][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N21
dffeas \my_reg[17][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][24] .is_wysiwyg = "true";
defparam \my_reg[17][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N20
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[25][24]~q )) # (!dcifimemload_24 & ((\my_reg[17][24]~q )))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[25][24]~q ),
	.datac(\my_reg[17][24]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hEE50;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N30
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// \Mux7~1_combout  = (dcifimemload_23 & ((\Mux7~0_combout  & ((\my_reg[29][24]~q ))) # (!\Mux7~0_combout  & (\my_reg[21][24]~q )))) # (!dcifimemload_23 & (((\Mux7~0_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[21][24]~q ),
	.datac(\my_reg[29][24]~q ),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hF588;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N13
dffeas \my_reg[23][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][24] .is_wysiwyg = "true";
defparam \my_reg[23][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N11
dffeas \my_reg[31][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][24] .is_wysiwyg = "true";
defparam \my_reg[31][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N13
dffeas \my_reg[19][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][24] .is_wysiwyg = "true";
defparam \my_reg[19][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N12
cycloneive_lcell_comb \Mux7~7 (
// Equation(s):
// \Mux7~7_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[27][24]~q )) # (!dcifimemload_24 & ((\my_reg[19][24]~q )))))

	.dataa(\my_reg[27][24]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[19][24]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux7~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~7 .lut_mask = 16'hEE30;
defparam \Mux7~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N10
cycloneive_lcell_comb \Mux7~8 (
// Equation(s):
// \Mux7~8_combout  = (dcifimemload_23 & ((\Mux7~7_combout  & ((\my_reg[31][24]~q ))) # (!\Mux7~7_combout  & (\my_reg[23][24]~q )))) # (!dcifimemload_23 & (((\Mux7~7_combout ))))

	.dataa(\my_reg[23][24]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[31][24]~q ),
	.datad(\Mux7~7_combout ),
	.cin(gnd),
	.combout(\Mux7~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~8 .lut_mask = 16'hF388;
defparam \Mux7~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N9
dffeas \my_reg[24][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][24] .is_wysiwyg = "true";
defparam \my_reg[24][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N11
dffeas \my_reg[28][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][24] .is_wysiwyg = "true";
defparam \my_reg[28][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N25
dffeas \my_reg[16][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][24] .is_wysiwyg = "true";
defparam \my_reg[16][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N24
cycloneive_lcell_comb \Mux7~4 (
// Equation(s):
// \Mux7~4_combout  = (dcifimemload_23 & ((\my_reg[20][24]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[16][24]~q  & !dcifimemload_24))))

	.dataa(\my_reg[20][24]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[16][24]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux7~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~4 .lut_mask = 16'hCCB8;
defparam \Mux7~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N10
cycloneive_lcell_comb \Mux7~5 (
// Equation(s):
// \Mux7~5_combout  = (dcifimemload_24 & ((\Mux7~4_combout  & ((\my_reg[28][24]~q ))) # (!\Mux7~4_combout  & (\my_reg[24][24]~q )))) # (!dcifimemload_24 & (((\Mux7~4_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[24][24]~q ),
	.datac(\my_reg[28][24]~q ),
	.datad(\Mux7~4_combout ),
	.cin(gnd),
	.combout(\Mux7~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~5 .lut_mask = 16'hF588;
defparam \Mux7~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N21
dffeas \my_reg[30][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][24] .is_wysiwyg = "true";
defparam \my_reg[30][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N3
dffeas \my_reg[18][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][24] .is_wysiwyg = "true";
defparam \my_reg[18][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N2
cycloneive_lcell_comb \Mux7~2 (
// Equation(s):
// \Mux7~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[22][24]~q )) # (!dcifimemload_23 & ((\my_reg[18][24]~q )))))

	.dataa(\my_reg[22][24]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[18][24]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~2 .lut_mask = 16'hEE30;
defparam \Mux7~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N20
cycloneive_lcell_comb \Mux7~3 (
// Equation(s):
// \Mux7~3_combout  = (dcifimemload_24 & ((\Mux7~2_combout  & ((\my_reg[30][24]~q ))) # (!\Mux7~2_combout  & (\my_reg[26][24]~q )))) # (!dcifimemload_24 & (((\Mux7~2_combout ))))

	.dataa(\my_reg[26][24]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[30][24]~q ),
	.datad(\Mux7~2_combout ),
	.cin(gnd),
	.combout(\Mux7~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~3 .lut_mask = 16'hF388;
defparam \Mux7~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N20
cycloneive_lcell_comb \Mux7~6 (
// Equation(s):
// \Mux7~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux7~3_combout ))) # (!dcifimemload_22 & (\Mux7~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux7~5_combout ),
	.datad(\Mux7~3_combout ),
	.cin(gnd),
	.combout(\Mux7~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~6 .lut_mask = 16'hDC98;
defparam \Mux7~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N11
dffeas \my_reg[7][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][24] .is_wysiwyg = "true";
defparam \my_reg[7][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N23
dffeas \my_reg[6][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][24] .is_wysiwyg = "true";
defparam \my_reg[6][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N1
dffeas \my_reg[4][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][24] .is_wysiwyg = "true";
defparam \my_reg[4][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N1
dffeas \my_reg[5][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][24] .is_wysiwyg = "true";
defparam \my_reg[5][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N0
cycloneive_lcell_comb \Mux7~10 (
// Equation(s):
// \Mux7~10_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\my_reg[5][24]~q ))) # (!dcifimemload_21 & (\my_reg[4][24]~q ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[4][24]~q ),
	.datac(\my_reg[5][24]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux7~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~10 .lut_mask = 16'hFA44;
defparam \Mux7~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N22
cycloneive_lcell_comb \Mux7~11 (
// Equation(s):
// \Mux7~11_combout  = (dcifimemload_22 & ((\Mux7~10_combout  & (\my_reg[7][24]~q )) # (!\Mux7~10_combout  & ((\my_reg[6][24]~q ))))) # (!dcifimemload_22 & (((\Mux7~10_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[7][24]~q ),
	.datac(\my_reg[6][24]~q ),
	.datad(\Mux7~10_combout ),
	.cin(gnd),
	.combout(\Mux7~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~11 .lut_mask = 16'hDDA0;
defparam \Mux7~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y31_N1
dffeas \my_reg[15][24] (
	.clk(CLK),
	.d(wdat9),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][24] .is_wysiwyg = "true";
defparam \my_reg[15][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N2
cycloneive_lcell_comb \my_reg[14][24]~feeder (
// Equation(s):
// \my_reg[14][24]~feeder_combout  = \wdat~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat9),
	.cin(gnd),
	.combout(\my_reg[14][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[14][24]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[14][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N3
dffeas \my_reg[14][24] (
	.clk(CLK),
	.d(\my_reg[14][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][24] .is_wysiwyg = "true";
defparam \my_reg[14][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N18
cycloneive_lcell_comb \my_reg[12][24]~feeder (
// Equation(s):
// \my_reg[12][24]~feeder_combout  = \wdat~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat9),
	.cin(gnd),
	.combout(\my_reg[12][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[12][24]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[12][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N19
dffeas \my_reg[12][24] (
	.clk(CLK),
	.d(\my_reg[12][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][24] .is_wysiwyg = "true";
defparam \my_reg[12][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N3
dffeas \my_reg[13][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][24] .is_wysiwyg = "true";
defparam \my_reg[13][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N16
cycloneive_lcell_comb \Mux7~17 (
// Equation(s):
// \Mux7~17_combout  = (dcifimemload_21 & (((\my_reg[13][24]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\my_reg[12][24]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[12][24]~q ),
	.datac(\my_reg[13][24]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux7~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~17 .lut_mask = 16'hAAE4;
defparam \Mux7~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N10
cycloneive_lcell_comb \Mux7~18 (
// Equation(s):
// \Mux7~18_combout  = (dcifimemload_22 & ((\Mux7~17_combout  & (\my_reg[15][24]~q )) # (!\Mux7~17_combout  & ((\my_reg[14][24]~q ))))) # (!dcifimemload_22 & (((\Mux7~17_combout ))))

	.dataa(\my_reg[15][24]~q ),
	.datab(\my_reg[14][24]~q ),
	.datac(dcifimemload_22),
	.datad(\Mux7~17_combout ),
	.cin(gnd),
	.combout(\Mux7~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~18 .lut_mask = 16'hAFC0;
defparam \Mux7~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y42_N7
dffeas \my_reg[9][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][24] .is_wysiwyg = "true";
defparam \my_reg[9][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y41_N23
dffeas \my_reg[11][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][24] .is_wysiwyg = "true";
defparam \my_reg[11][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y42_N9
dffeas \my_reg[10][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][24] .is_wysiwyg = "true";
defparam \my_reg[10][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y41_N1
dffeas \my_reg[8][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][24] .is_wysiwyg = "true";
defparam \my_reg[8][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N0
cycloneive_lcell_comb \Mux7~12 (
// Equation(s):
// \Mux7~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][24]~q )) # (!dcifimemload_22 & ((\my_reg[8][24]~q )))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[10][24]~q ),
	.datac(\my_reg[8][24]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux7~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~12 .lut_mask = 16'hEE50;
defparam \Mux7~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N22
cycloneive_lcell_comb \Mux7~13 (
// Equation(s):
// \Mux7~13_combout  = (dcifimemload_21 & ((\Mux7~12_combout  & ((\my_reg[11][24]~q ))) # (!\Mux7~12_combout  & (\my_reg[9][24]~q )))) # (!dcifimemload_21 & (((\Mux7~12_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][24]~q ),
	.datac(\my_reg[11][24]~q ),
	.datad(\Mux7~12_combout ),
	.cin(gnd),
	.combout(\Mux7~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~13 .lut_mask = 16'hF588;
defparam \Mux7~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N15
dffeas \my_reg[2][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][24] .is_wysiwyg = "true";
defparam \my_reg[2][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N23
dffeas \my_reg[1][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][24] .is_wysiwyg = "true";
defparam \my_reg[1][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N22
cycloneive_lcell_comb \Mux7~14 (
// Equation(s):
// \Mux7~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\my_reg[3][24]~q )) # (!dcifimemload_22 & ((\my_reg[1][24]~q )))))

	.dataa(\my_reg[3][24]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[1][24]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux7~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~14 .lut_mask = 16'h88C0;
defparam \Mux7~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N14
cycloneive_lcell_comb \Mux7~15 (
// Equation(s):
// \Mux7~15_combout  = (\Mux7~14_combout ) # ((dcifimemload_22 & (!dcifimemload_21 & \my_reg[2][24]~q )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\my_reg[2][24]~q ),
	.datad(\Mux7~14_combout ),
	.cin(gnd),
	.combout(\Mux7~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~15 .lut_mask = 16'hFF20;
defparam \Mux7~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N12
cycloneive_lcell_comb \Mux7~16 (
// Equation(s):
// \Mux7~16_combout  = (dcifimemload_23 & (dcifimemload_24)) # (!dcifimemload_23 & ((dcifimemload_24 & (\Mux7~13_combout )) # (!dcifimemload_24 & ((\Mux7~15_combout )))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux7~13_combout ),
	.datad(\Mux7~15_combout ),
	.cin(gnd),
	.combout(\Mux7~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~16 .lut_mask = 16'hD9C8;
defparam \Mux7~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N17
dffeas \my_reg[3][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][24] .is_wysiwyg = "true";
defparam \my_reg[3][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N16
cycloneive_lcell_comb \Mux39~4 (
// Equation(s):
// \Mux39~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][24]~q ))) # (!dcifimemload_17 & (\my_reg[1][24]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[1][24]~q ),
	.datac(\my_reg[3][24]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux39~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~4 .lut_mask = 16'hE400;
defparam \Mux39~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N8
cycloneive_lcell_comb \Mux39~5 (
// Equation(s):
// \Mux39~5_combout  = (\Mux39~4_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \my_reg[2][24]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux39~4_combout ),
	.datad(\my_reg[2][24]~q ),
	.cin(gnd),
	.combout(\Mux39~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~5 .lut_mask = 16'hF2F0;
defparam \Mux39~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N0
cycloneive_lcell_comb \Mux39~2 (
// Equation(s):
// \Mux39~2_combout  = (dcifimemload_16 & ((\my_reg[5][24]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\my_reg[4][24]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[5][24]~q ),
	.datac(\my_reg[4][24]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux39~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~2 .lut_mask = 16'hAAD8;
defparam \Mux39~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N10
cycloneive_lcell_comb \Mux39~3 (
// Equation(s):
// \Mux39~3_combout  = (dcifimemload_17 & ((\Mux39~2_combout  & ((\my_reg[7][24]~q ))) # (!\Mux39~2_combout  & (\my_reg[6][24]~q )))) # (!dcifimemload_17 & (((\Mux39~2_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[6][24]~q ),
	.datac(\my_reg[7][24]~q ),
	.datad(\Mux39~2_combout ),
	.cin(gnd),
	.combout(\Mux39~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~3 .lut_mask = 16'hF588;
defparam \Mux39~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N30
cycloneive_lcell_comb \Mux39~6 (
// Equation(s):
// \Mux39~6_combout  = (dcifimemload_18 & ((dcifimemload_19) # ((\Mux39~3_combout )))) # (!dcifimemload_18 & (!dcifimemload_19 & (\Mux39~5_combout )))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux39~5_combout ),
	.datad(\Mux39~3_combout ),
	.cin(gnd),
	.combout(\Mux39~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~6 .lut_mask = 16'hBA98;
defparam \Mux39~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N2
cycloneive_lcell_comb \Mux39~7 (
// Equation(s):
// \Mux39~7_combout  = (dcifimemload_16 & (((\my_reg[13][24]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[12][24]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[12][24]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[13][24]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux39~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~7 .lut_mask = 16'hCCE2;
defparam \Mux39~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N6
cycloneive_lcell_comb \Mux39~8 (
// Equation(s):
// \Mux39~8_combout  = (dcifimemload_17 & ((\Mux39~7_combout  & (\my_reg[15][24]~q )) # (!\Mux39~7_combout  & ((\my_reg[14][24]~q ))))) # (!dcifimemload_17 & (((\Mux39~7_combout ))))

	.dataa(\my_reg[15][24]~q ),
	.datab(\my_reg[14][24]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux39~7_combout ),
	.cin(gnd),
	.combout(\Mux39~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~8 .lut_mask = 16'hAFC0;
defparam \Mux39~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N8
cycloneive_lcell_comb \Mux39~0 (
// Equation(s):
// \Mux39~0_combout  = (dcifimemload_17 & (((\my_reg[10][24]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\my_reg[8][24]~q  & ((!dcifimemload_16))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[8][24]~q ),
	.datac(\my_reg[10][24]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux39~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~0 .lut_mask = 16'hAAE4;
defparam \Mux39~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N6
cycloneive_lcell_comb \Mux39~1 (
// Equation(s):
// \Mux39~1_combout  = (\Mux39~0_combout  & ((\my_reg[11][24]~q ) # ((!dcifimemload_16)))) # (!\Mux39~0_combout  & (((\my_reg[9][24]~q  & dcifimemload_16))))

	.dataa(\my_reg[11][24]~q ),
	.datab(\Mux39~0_combout ),
	.datac(\my_reg[9][24]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux39~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~1 .lut_mask = 16'hB8CC;
defparam \Mux39~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N0
cycloneive_lcell_comb \Mux39~10 (
// Equation(s):
// \Mux39~10_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[21][24]~q ))) # (!dcifimemload_18 & (\my_reg[17][24]~q ))))

	.dataa(\my_reg[17][24]~q ),
	.datab(\my_reg[21][24]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux39~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~10 .lut_mask = 16'hFC0A;
defparam \Mux39~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N0
cycloneive_lcell_comb \Mux39~11 (
// Equation(s):
// \Mux39~11_combout  = (\Mux39~10_combout  & ((\my_reg[29][24]~q ) # ((!dcifimemload_19)))) # (!\Mux39~10_combout  & (((\my_reg[25][24]~q  & dcifimemload_19))))

	.dataa(\my_reg[29][24]~q ),
	.datab(\my_reg[25][24]~q ),
	.datac(\Mux39~10_combout ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux39~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~11 .lut_mask = 16'hACF0;
defparam \Mux39~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N23
dffeas \my_reg[27][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][24] .is_wysiwyg = "true";
defparam \my_reg[27][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N12
cycloneive_lcell_comb \Mux39~17 (
// Equation(s):
// \Mux39~17_combout  = (dcifimemload_18 & (((\my_reg[23][24]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[19][24]~q  & ((!dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[19][24]~q ),
	.datac(\my_reg[23][24]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux39~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~17 .lut_mask = 16'hAAE4;
defparam \Mux39~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N22
cycloneive_lcell_comb \Mux39~18 (
// Equation(s):
// \Mux39~18_combout  = (dcifimemload_19 & ((\Mux39~17_combout  & (\my_reg[31][24]~q )) # (!\Mux39~17_combout  & ((\my_reg[27][24]~q ))))) # (!dcifimemload_19 & (((\Mux39~17_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[31][24]~q ),
	.datac(\my_reg[27][24]~q ),
	.datad(\Mux39~17_combout ),
	.cin(gnd),
	.combout(\Mux39~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~18 .lut_mask = 16'hDDA0;
defparam \Mux39~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N8
cycloneive_lcell_comb \Mux39~14 (
// Equation(s):
// \Mux39~14_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & (\my_reg[24][24]~q )) # (!dcifimemload_19 & ((\my_reg[16][24]~q )))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\my_reg[24][24]~q ),
	.datad(\my_reg[16][24]~q ),
	.cin(gnd),
	.combout(\Mux39~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~14 .lut_mask = 16'hD9C8;
defparam \Mux39~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N15
dffeas \my_reg[20][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][24] .is_wysiwyg = "true";
defparam \my_reg[20][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N14
cycloneive_lcell_comb \Mux39~15 (
// Equation(s):
// \Mux39~15_combout  = (\Mux39~14_combout  & ((\my_reg[28][24]~q ) # ((!dcifimemload_18)))) # (!\Mux39~14_combout  & (((\my_reg[20][24]~q  & dcifimemload_18))))

	.dataa(\my_reg[28][24]~q ),
	.datab(\Mux39~14_combout ),
	.datac(\my_reg[20][24]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux39~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~15 .lut_mask = 16'hB8CC;
defparam \Mux39~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N23
dffeas \my_reg[22][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][24] .is_wysiwyg = "true";
defparam \my_reg[22][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N5
dffeas \my_reg[26][24] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][24] .is_wysiwyg = "true";
defparam \my_reg[26][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N4
cycloneive_lcell_comb \Mux39~12 (
// Equation(s):
// \Mux39~12_combout  = (dcifimemload_19 & (((\my_reg[26][24]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[18][24]~q  & ((!dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[18][24]~q ),
	.datac(\my_reg[26][24]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux39~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~12 .lut_mask = 16'hAAE4;
defparam \Mux39~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N22
cycloneive_lcell_comb \Mux39~13 (
// Equation(s):
// \Mux39~13_combout  = (dcifimemload_18 & ((\Mux39~12_combout  & (\my_reg[30][24]~q )) # (!\Mux39~12_combout  & ((\my_reg[22][24]~q ))))) # (!dcifimemload_18 & (((\Mux39~12_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[30][24]~q ),
	.datac(\my_reg[22][24]~q ),
	.datad(\Mux39~12_combout ),
	.cin(gnd),
	.combout(\Mux39~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~13 .lut_mask = 16'hDDA0;
defparam \Mux39~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N16
cycloneive_lcell_comb \Mux39~16 (
// Equation(s):
// \Mux39~16_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux39~13_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & (\Mux39~15_combout )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux39~15_combout ),
	.datad(\Mux39~13_combout ),
	.cin(gnd),
	.combout(\Mux39~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~16 .lut_mask = 16'hBA98;
defparam \Mux39~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N11
dffeas \my_reg[11][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][23] .is_wysiwyg = "true";
defparam \my_reg[11][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N8
cycloneive_lcell_comb \my_reg[9][23]~feeder (
// Equation(s):
// \my_reg[9][23]~feeder_combout  = \wdat~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat10),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[9][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[9][23]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[9][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N9
dffeas \my_reg[9][23] (
	.clk(CLK),
	.d(\my_reg[9][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][23] .is_wysiwyg = "true";
defparam \my_reg[9][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N10
cycloneive_lcell_comb \Mux8~11 (
// Equation(s):
// \Mux8~11_combout  = (\Mux8~10_combout  & ((\my_reg[11][23]~q ) # ((!dcifimemload_21)))) # (!\Mux8~10_combout  & (((dcifimemload_21 & \my_reg[9][23]~q ))))

	.dataa(\Mux8~10_combout ),
	.datab(\my_reg[11][23]~q ),
	.datac(dcifimemload_21),
	.datad(\my_reg[9][23]~q ),
	.cin(gnd),
	.combout(\Mux8~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~11 .lut_mask = 16'hDA8A;
defparam \Mux8~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N25
dffeas \my_reg[14][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][23] .is_wysiwyg = "true";
defparam \my_reg[14][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N31
dffeas \my_reg[15][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][23] .is_wysiwyg = "true";
defparam \my_reg[15][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N20
cycloneive_lcell_comb \my_reg[12][23]~feeder (
// Equation(s):
// \my_reg[12][23]~feeder_combout  = \wdat~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat10),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[12][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[12][23]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[12][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N21
dffeas \my_reg[12][23] (
	.clk(CLK),
	.d(\my_reg[12][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][23] .is_wysiwyg = "true";
defparam \my_reg[12][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N14
cycloneive_lcell_comb \Mux8~17 (
// Equation(s):
// \Mux8~17_combout  = (dcifimemload_21 & ((\my_reg[13][23]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][23]~q  & !dcifimemload_22))))

	.dataa(\my_reg[13][23]~q ),
	.datab(\my_reg[12][23]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux8~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~17 .lut_mask = 16'hF0AC;
defparam \Mux8~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N30
cycloneive_lcell_comb \Mux8~18 (
// Equation(s):
// \Mux8~18_combout  = (dcifimemload_22 & ((\Mux8~17_combout  & ((\my_reg[15][23]~q ))) # (!\Mux8~17_combout  & (\my_reg[14][23]~q )))) # (!dcifimemload_22 & (((\Mux8~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[14][23]~q ),
	.datac(\my_reg[15][23]~q ),
	.datad(\Mux8~17_combout ),
	.cin(gnd),
	.combout(\Mux8~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~18 .lut_mask = 16'hF588;
defparam \Mux8~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N5
dffeas \my_reg[6][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][23] .is_wysiwyg = "true";
defparam \my_reg[6][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N13
dffeas \my_reg[7][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][23] .is_wysiwyg = "true";
defparam \my_reg[7][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N4
cycloneive_lcell_comb \my_reg[4][23]~feeder (
// Equation(s):
// \my_reg[4][23]~feeder_combout  = \wdat~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat10),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[4][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[4][23]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[4][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y42_N5
dffeas \my_reg[4][23] (
	.clk(CLK),
	.d(\my_reg[4][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][23] .is_wysiwyg = "true";
defparam \my_reg[4][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N6
cycloneive_lcell_comb \Mux8~12 (
// Equation(s):
// \Mux8~12_combout  = (dcifimemload_21 & ((\my_reg[5][23]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[4][23]~q  & !dcifimemload_22))))

	.dataa(\my_reg[5][23]~q ),
	.datab(\my_reg[4][23]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux8~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~12 .lut_mask = 16'hF0AC;
defparam \Mux8~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N12
cycloneive_lcell_comb \Mux8~13 (
// Equation(s):
// \Mux8~13_combout  = (dcifimemload_22 & ((\Mux8~12_combout  & ((\my_reg[7][23]~q ))) # (!\Mux8~12_combout  & (\my_reg[6][23]~q )))) # (!dcifimemload_22 & (((\Mux8~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[6][23]~q ),
	.datac(\my_reg[7][23]~q ),
	.datad(\Mux8~12_combout ),
	.cin(gnd),
	.combout(\Mux8~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~13 .lut_mask = 16'hF588;
defparam \Mux8~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N29
dffeas \my_reg[3][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][23] .is_wysiwyg = "true";
defparam \my_reg[3][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N25
dffeas \my_reg[1][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][23] .is_wysiwyg = "true";
defparam \my_reg[1][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N24
cycloneive_lcell_comb \Mux8~14 (
// Equation(s):
// \Mux8~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\my_reg[3][23]~q )) # (!dcifimemload_22 & ((\my_reg[1][23]~q )))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[3][23]~q ),
	.datac(\my_reg[1][23]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux8~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~14 .lut_mask = 16'h88A0;
defparam \Mux8~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y39_N19
dffeas \my_reg[2][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][23] .is_wysiwyg = "true";
defparam \my_reg[2][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N18
cycloneive_lcell_comb \Mux8~15 (
// Equation(s):
// \Mux8~15_combout  = (\Mux8~14_combout ) # ((!dcifimemload_21 & (\my_reg[2][23]~q  & dcifimemload_22)))

	.dataa(dcifimemload_21),
	.datab(\Mux8~14_combout ),
	.datac(\my_reg[2][23]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux8~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~15 .lut_mask = 16'hDCCC;
defparam \Mux8~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N0
cycloneive_lcell_comb \Mux8~16 (
// Equation(s):
// \Mux8~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & (\Mux8~13_combout )) # (!dcifimemload_23 & ((\Mux8~15_combout )))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux8~13_combout ),
	.datad(\Mux8~15_combout ),
	.cin(gnd),
	.combout(\Mux8~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~16 .lut_mask = 16'hD9C8;
defparam \Mux8~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N2
cycloneive_lcell_comb \Mux8~19 (
// Equation(s):
// \Mux8~19_combout  = (dcifimemload_24 & ((\Mux8~16_combout  & ((\Mux8~18_combout ))) # (!\Mux8~16_combout  & (\Mux8~11_combout )))) # (!dcifimemload_24 & (((\Mux8~16_combout ))))

	.dataa(dcifimemload_24),
	.datab(\Mux8~11_combout ),
	.datac(\Mux8~18_combout ),
	.datad(\Mux8~16_combout ),
	.cin(gnd),
	.combout(\Mux8~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~19 .lut_mask = 16'hF588;
defparam \Mux8~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N1
dffeas \my_reg[27][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][23] .is_wysiwyg = "true";
defparam \my_reg[27][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y41_N11
dffeas \my_reg[31][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][23] .is_wysiwyg = "true";
defparam \my_reg[31][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N11
dffeas \my_reg[23][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][23] .is_wysiwyg = "true";
defparam \my_reg[23][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y41_N21
dffeas \my_reg[19][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][23] .is_wysiwyg = "true";
defparam \my_reg[19][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N20
cycloneive_lcell_comb \Mux8~7 (
// Equation(s):
// \Mux8~7_combout  = (dcifimemload_23 & ((\my_reg[23][23]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[19][23]~q  & !dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[23][23]~q ),
	.datac(\my_reg[19][23]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux8~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~7 .lut_mask = 16'hAAD8;
defparam \Mux8~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N10
cycloneive_lcell_comb \Mux8~8 (
// Equation(s):
// \Mux8~8_combout  = (dcifimemload_24 & ((\Mux8~7_combout  & ((\my_reg[31][23]~q ))) # (!\Mux8~7_combout  & (\my_reg[27][23]~q )))) # (!dcifimemload_24 & (((\Mux8~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[27][23]~q ),
	.datac(\my_reg[31][23]~q ),
	.datad(\Mux8~7_combout ),
	.cin(gnd),
	.combout(\Mux8~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~8 .lut_mask = 16'hF588;
defparam \Mux8~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N28
cycloneive_lcell_comb \my_reg[25][23]~feeder (
// Equation(s):
// \my_reg[25][23]~feeder_combout  = \wdat~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat10),
	.cin(gnd),
	.combout(\my_reg[25][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][23]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[25][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N29
dffeas \my_reg[25][23] (
	.clk(CLK),
	.d(\my_reg[25][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][23] .is_wysiwyg = "true";
defparam \my_reg[25][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N17
dffeas \my_reg[29][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][23] .is_wysiwyg = "true";
defparam \my_reg[29][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N19
dffeas \my_reg[17][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][23] .is_wysiwyg = "true";
defparam \my_reg[17][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N18
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (dcifimemload_23 & ((\my_reg[21][23]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[17][23]~q  & !dcifimemload_24))))

	.dataa(\my_reg[21][23]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[17][23]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hCCB8;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N16
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// \Mux8~1_combout  = (dcifimemload_24 & ((\Mux8~0_combout  & ((\my_reg[29][23]~q ))) # (!\Mux8~0_combout  & (\my_reg[25][23]~q )))) # (!dcifimemload_24 & (((\Mux8~0_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[25][23]~q ),
	.datac(\my_reg[29][23]~q ),
	.datad(\Mux8~0_combout ),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hF588;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y30_N31
dffeas \my_reg[28][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][23] .is_wysiwyg = "true";
defparam \my_reg[28][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N17
dffeas \my_reg[16][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][23] .is_wysiwyg = "true";
defparam \my_reg[16][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N16
cycloneive_lcell_comb \Mux8~4 (
// Equation(s):
// \Mux8~4_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[24][23]~q )) # (!dcifimemload_24 & ((\my_reg[16][23]~q )))))

	.dataa(\my_reg[24][23]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[16][23]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~4 .lut_mask = 16'hEE30;
defparam \Mux8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N30
cycloneive_lcell_comb \Mux8~5 (
// Equation(s):
// \Mux8~5_combout  = (dcifimemload_23 & ((\Mux8~4_combout  & ((\my_reg[28][23]~q ))) # (!\Mux8~4_combout  & (\my_reg[20][23]~q )))) # (!dcifimemload_23 & (((\Mux8~4_combout ))))

	.dataa(\my_reg[20][23]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[28][23]~q ),
	.datad(\Mux8~4_combout ),
	.cin(gnd),
	.combout(\Mux8~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~5 .lut_mask = 16'hF388;
defparam \Mux8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y42_N25
dffeas \my_reg[22][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][23] .is_wysiwyg = "true";
defparam \my_reg[22][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N11
dffeas \my_reg[30][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][23] .is_wysiwyg = "true";
defparam \my_reg[30][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y42_N7
dffeas \my_reg[26][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][23] .is_wysiwyg = "true";
defparam \my_reg[26][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N21
dffeas \my_reg[18][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][23] .is_wysiwyg = "true";
defparam \my_reg[18][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N20
cycloneive_lcell_comb \Mux8~2 (
// Equation(s):
// \Mux8~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[26][23]~q )) # (!dcifimemload_24 & ((\my_reg[18][23]~q )))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[26][23]~q ),
	.datac(\my_reg[18][23]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux8~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~2 .lut_mask = 16'hEE50;
defparam \Mux8~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N10
cycloneive_lcell_comb \Mux8~3 (
// Equation(s):
// \Mux8~3_combout  = (dcifimemload_23 & ((\Mux8~2_combout  & ((\my_reg[30][23]~q ))) # (!\Mux8~2_combout  & (\my_reg[22][23]~q )))) # (!dcifimemload_23 & (((\Mux8~2_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[22][23]~q ),
	.datac(\my_reg[30][23]~q ),
	.datad(\Mux8~2_combout ),
	.cin(gnd),
	.combout(\Mux8~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~3 .lut_mask = 16'hF588;
defparam \Mux8~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N2
cycloneive_lcell_comb \Mux8~6 (
// Equation(s):
// \Mux8~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux8~3_combout ))) # (!dcifimemload_22 & (\Mux8~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux8~5_combout ),
	.datad(\Mux8~3_combout ),
	.cin(gnd),
	.combout(\Mux8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~6 .lut_mask = 16'hDC98;
defparam \Mux8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N24
cycloneive_lcell_comb \Mux8~9 (
// Equation(s):
// \Mux8~9_combout  = (dcifimemload_21 & ((\Mux8~6_combout  & (\Mux8~8_combout )) # (!\Mux8~6_combout  & ((\Mux8~1_combout ))))) # (!dcifimemload_21 & (((\Mux8~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux8~8_combout ),
	.datac(\Mux8~1_combout ),
	.datad(\Mux8~6_combout ),
	.cin(gnd),
	.combout(\Mux8~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~9 .lut_mask = 16'hDDA0;
defparam \Mux8~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N19
dffeas \my_reg[5][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][23] .is_wysiwyg = "true";
defparam \my_reg[5][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N18
cycloneive_lcell_comb \Mux40~0 (
// Equation(s):
// \Mux40~0_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][23]~q ))) # (!dcifimemload_16 & (\my_reg[4][23]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[4][23]~q ),
	.datac(\my_reg[5][23]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux40~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~0 .lut_mask = 16'hFA44;
defparam \Mux40~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N4
cycloneive_lcell_comb \Mux40~1 (
// Equation(s):
// \Mux40~1_combout  = (dcifimemload_17 & ((\Mux40~0_combout  & (\my_reg[7][23]~q )) # (!\Mux40~0_combout  & ((\my_reg[6][23]~q ))))) # (!dcifimemload_17 & (((\Mux40~0_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[7][23]~q ),
	.datac(\my_reg[6][23]~q ),
	.datad(\Mux40~0_combout ),
	.cin(gnd),
	.combout(\Mux40~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~1 .lut_mask = 16'hDDA0;
defparam \Mux40~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N4
cycloneive_lcell_comb \my_reg[10][23]~feeder (
// Equation(s):
// \my_reg[10][23]~feeder_combout  = \wdat~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat10),
	.cin(gnd),
	.combout(\my_reg[10][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[10][23]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[10][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y38_N5
dffeas \my_reg[10][23] (
	.clk(CLK),
	.d(\my_reg[10][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][23] .is_wysiwyg = "true";
defparam \my_reg[10][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N17
dffeas \my_reg[8][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][23] .is_wysiwyg = "true";
defparam \my_reg[8][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N16
cycloneive_lcell_comb \Mux40~2 (
// Equation(s):
// \Mux40~2_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\my_reg[10][23]~q )) # (!dcifimemload_17 & ((\my_reg[8][23]~q )))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[10][23]~q ),
	.datac(\my_reg[8][23]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux40~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~2 .lut_mask = 16'hEE50;
defparam \Mux40~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N10
cycloneive_lcell_comb \Mux40~3 (
// Equation(s):
// \Mux40~3_combout  = (\Mux40~2_combout  & (((\my_reg[11][23]~q ) # (!dcifimemload_16)))) # (!\Mux40~2_combout  & (\my_reg[9][23]~q  & ((dcifimemload_16))))

	.dataa(\my_reg[9][23]~q ),
	.datab(\Mux40~2_combout ),
	.datac(\my_reg[11][23]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux40~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~3 .lut_mask = 16'hE2CC;
defparam \Mux40~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N28
cycloneive_lcell_comb \Mux40~4 (
// Equation(s):
// \Mux40~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][23]~q ))) # (!dcifimemload_17 & (\my_reg[1][23]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[1][23]~q ),
	.datac(\my_reg[3][23]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux40~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~4 .lut_mask = 16'hE400;
defparam \Mux40~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N2
cycloneive_lcell_comb \Mux40~5 (
// Equation(s):
// \Mux40~5_combout  = (\Mux40~4_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \my_reg[2][23]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux40~4_combout ),
	.datad(\my_reg[2][23]~q ),
	.cin(gnd),
	.combout(\Mux40~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~5 .lut_mask = 16'hF2F0;
defparam \Mux40~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N4
cycloneive_lcell_comb \Mux40~6 (
// Equation(s):
// \Mux40~6_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & (\Mux40~3_combout )) # (!dcifimemload_19 & ((\Mux40~5_combout )))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux40~3_combout ),
	.datad(\Mux40~5_combout ),
	.cin(gnd),
	.combout(\Mux40~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~6 .lut_mask = 16'hD9C8;
defparam \Mux40~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N24
cycloneive_lcell_comb \Mux40~7 (
// Equation(s):
// \Mux40~7_combout  = (dcifimemload_16 & ((\my_reg[13][23]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\my_reg[12][23]~q  & !dcifimemload_17))))

	.dataa(\my_reg[13][23]~q ),
	.datab(\my_reg[12][23]~q ),
	.datac(dcifimemload_16),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux40~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~7 .lut_mask = 16'hF0AC;
defparam \Mux40~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N24
cycloneive_lcell_comb \Mux40~8 (
// Equation(s):
// \Mux40~8_combout  = (dcifimemload_17 & ((\Mux40~7_combout  & (\my_reg[15][23]~q )) # (!\Mux40~7_combout  & ((\my_reg[14][23]~q ))))) # (!dcifimemload_17 & (((\Mux40~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[15][23]~q ),
	.datac(\my_reg[14][23]~q ),
	.datad(\Mux40~7_combout ),
	.cin(gnd),
	.combout(\Mux40~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~8 .lut_mask = 16'hDDA0;
defparam \Mux40~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N0
cycloneive_lcell_comb \Mux40~17 (
// Equation(s):
// \Mux40~17_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[27][23]~q ))) # (!dcifimemload_19 & (\my_reg[19][23]~q ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[19][23]~q ),
	.datac(\my_reg[27][23]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux40~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~17 .lut_mask = 16'hFA44;
defparam \Mux40~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N10
cycloneive_lcell_comb \Mux40~18 (
// Equation(s):
// \Mux40~18_combout  = (dcifimemload_18 & ((\Mux40~17_combout  & (\my_reg[31][23]~q )) # (!\Mux40~17_combout  & ((\my_reg[23][23]~q ))))) # (!dcifimemload_18 & (((\Mux40~17_combout ))))

	.dataa(\my_reg[31][23]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[23][23]~q ),
	.datad(\Mux40~17_combout ),
	.cin(gnd),
	.combout(\Mux40~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~18 .lut_mask = 16'hBBC0;
defparam \Mux40~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N22
cycloneive_lcell_comb \Mux40~10 (
// Equation(s):
// \Mux40~10_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\my_reg[25][23]~q )) # (!dcifimemload_19 & ((\my_reg[17][23]~q )))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[25][23]~q ),
	.datac(\my_reg[17][23]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux40~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~10 .lut_mask = 16'hEE50;
defparam \Mux40~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N11
dffeas \my_reg[21][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][23] .is_wysiwyg = "true";
defparam \my_reg[21][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N10
cycloneive_lcell_comb \Mux40~11 (
// Equation(s):
// \Mux40~11_combout  = (\Mux40~10_combout  & ((\my_reg[29][23]~q ) # ((!dcifimemload_18)))) # (!\Mux40~10_combout  & (((\my_reg[21][23]~q  & dcifimemload_18))))

	.dataa(\Mux40~10_combout ),
	.datab(\my_reg[29][23]~q ),
	.datac(\my_reg[21][23]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux40~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~11 .lut_mask = 16'hD8AA;
defparam \Mux40~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N11
dffeas \my_reg[24][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][23] .is_wysiwyg = "true";
defparam \my_reg[24][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y42_N29
dffeas \my_reg[20][23] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][23] .is_wysiwyg = "true";
defparam \my_reg[20][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N28
cycloneive_lcell_comb \Mux40~14 (
// Equation(s):
// \Mux40~14_combout  = (dcifimemload_18 & ((dcifimemload_19) # ((\my_reg[20][23]~q )))) # (!dcifimemload_18 & (!dcifimemload_19 & ((\my_reg[16][23]~q ))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\my_reg[20][23]~q ),
	.datad(\my_reg[16][23]~q ),
	.cin(gnd),
	.combout(\Mux40~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~14 .lut_mask = 16'hB9A8;
defparam \Mux40~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N10
cycloneive_lcell_comb \Mux40~15 (
// Equation(s):
// \Mux40~15_combout  = (dcifimemload_19 & ((\Mux40~14_combout  & (\my_reg[28][23]~q )) # (!\Mux40~14_combout  & ((\my_reg[24][23]~q ))))) # (!dcifimemload_19 & (((\Mux40~14_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[28][23]~q ),
	.datac(\my_reg[24][23]~q ),
	.datad(\Mux40~14_combout ),
	.cin(gnd),
	.combout(\Mux40~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~15 .lut_mask = 16'hDDA0;
defparam \Mux40~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N24
cycloneive_lcell_comb \Mux40~12 (
// Equation(s):
// \Mux40~12_combout  = (dcifimemload_18 & (((\my_reg[22][23]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[18][23]~q  & ((!dcifimemload_19))))

	.dataa(\my_reg[18][23]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[22][23]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux40~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~12 .lut_mask = 16'hCCE2;
defparam \Mux40~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N6
cycloneive_lcell_comb \Mux40~13 (
// Equation(s):
// \Mux40~13_combout  = (dcifimemload_19 & ((\Mux40~12_combout  & (\my_reg[30][23]~q )) # (!\Mux40~12_combout  & ((\my_reg[26][23]~q ))))) # (!dcifimemload_19 & (((\Mux40~12_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[30][23]~q ),
	.datac(\my_reg[26][23]~q ),
	.datad(\Mux40~12_combout ),
	.cin(gnd),
	.combout(\Mux40~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~13 .lut_mask = 16'hDDA0;
defparam \Mux40~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N24
cycloneive_lcell_comb \Mux40~16 (
// Equation(s):
// \Mux40~16_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux40~13_combout ))) # (!dcifimemload_17 & (\Mux40~15_combout ))))

	.dataa(\Mux40~15_combout ),
	.datab(dcifimemload_16),
	.datac(dcifimemload_17),
	.datad(\Mux40~13_combout ),
	.cin(gnd),
	.combout(\Mux40~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~16 .lut_mask = 16'hF2C2;
defparam \Mux40~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N18
cycloneive_lcell_comb \my_reg[15][22]~feeder (
// Equation(s):
// \my_reg[15][22]~feeder_combout  = \wdat~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat11),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[15][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[15][22]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[15][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N19
dffeas \my_reg[15][22] (
	.clk(CLK),
	.d(\my_reg[15][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][22] .is_wysiwyg = "true";
defparam \my_reg[15][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N31
dffeas \my_reg[13][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][22] .is_wysiwyg = "true";
defparam \my_reg[13][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N9
dffeas \my_reg[12][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][22] .is_wysiwyg = "true";
defparam \my_reg[12][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N8
cycloneive_lcell_comb \Mux9~17 (
// Equation(s):
// \Mux9~17_combout  = (dcifimemload_21 & ((\my_reg[13][22]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][22]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[13][22]~q ),
	.datac(\my_reg[12][22]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux9~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~17 .lut_mask = 16'hAAD8;
defparam \Mux9~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N22
cycloneive_lcell_comb \Mux9~18 (
// Equation(s):
// \Mux9~18_combout  = (\Mux9~17_combout  & (((\my_reg[15][22]~q ) # (!dcifimemload_22)))) # (!\Mux9~17_combout  & (\my_reg[14][22]~q  & ((dcifimemload_22))))

	.dataa(\my_reg[14][22]~q ),
	.datab(\my_reg[15][22]~q ),
	.datac(\Mux9~17_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux9~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~18 .lut_mask = 16'hCAF0;
defparam \Mux9~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N17
dffeas \my_reg[6][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][22] .is_wysiwyg = "true";
defparam \my_reg[6][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y43_N31
dffeas \my_reg[7][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][22] .is_wysiwyg = "true";
defparam \my_reg[7][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y43_N25
dffeas \my_reg[4][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][22] .is_wysiwyg = "true";
defparam \my_reg[4][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N24
cycloneive_lcell_comb \Mux9~10 (
// Equation(s):
// \Mux9~10_combout  = (dcifimemload_21 & ((\my_reg[5][22]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[4][22]~q  & !dcifimemload_22))))

	.dataa(\my_reg[5][22]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[4][22]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux9~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~10 .lut_mask = 16'hCCB8;
defparam \Mux9~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N30
cycloneive_lcell_comb \Mux9~11 (
// Equation(s):
// \Mux9~11_combout  = (dcifimemload_22 & ((\Mux9~10_combout  & ((\my_reg[7][22]~q ))) # (!\Mux9~10_combout  & (\my_reg[6][22]~q )))) # (!dcifimemload_22 & (((\Mux9~10_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[6][22]~q ),
	.datac(\my_reg[7][22]~q ),
	.datad(\Mux9~10_combout ),
	.cin(gnd),
	.combout(\Mux9~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~11 .lut_mask = 16'hF588;
defparam \Mux9~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N1
dffeas \my_reg[2][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][22] .is_wysiwyg = "true";
defparam \my_reg[2][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N5
dffeas \my_reg[1][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][22] .is_wysiwyg = "true";
defparam \my_reg[1][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N4
cycloneive_lcell_comb \Mux9~14 (
// Equation(s):
// \Mux9~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\my_reg[3][22]~q )) # (!dcifimemload_22 & ((\my_reg[1][22]~q )))))

	.dataa(\my_reg[3][22]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[1][22]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux9~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~14 .lut_mask = 16'h88C0;
defparam \Mux9~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N0
cycloneive_lcell_comb \Mux9~15 (
// Equation(s):
// \Mux9~15_combout  = (\Mux9~14_combout ) # ((!dcifimemload_21 & (dcifimemload_22 & \my_reg[2][22]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\my_reg[2][22]~q ),
	.datad(\Mux9~14_combout ),
	.cin(gnd),
	.combout(\Mux9~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~15 .lut_mask = 16'hFF40;
defparam \Mux9~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y42_N31
dffeas \my_reg[9][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][22] .is_wysiwyg = "true";
defparam \my_reg[9][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y41_N9
dffeas \my_reg[11][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][22] .is_wysiwyg = "true";
defparam \my_reg[11][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N0
cycloneive_lcell_comb \my_reg[10][22]~feeder (
// Equation(s):
// \my_reg[10][22]~feeder_combout  = \wdat~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat11),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[10][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[10][22]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[10][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y42_N1
dffeas \my_reg[10][22] (
	.clk(CLK),
	.d(\my_reg[10][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][22] .is_wysiwyg = "true";
defparam \my_reg[10][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y41_N19
dffeas \my_reg[8][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][22] .is_wysiwyg = "true";
defparam \my_reg[8][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N18
cycloneive_lcell_comb \Mux9~12 (
// Equation(s):
// \Mux9~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][22]~q )) # (!dcifimemload_22 & ((\my_reg[8][22]~q )))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[10][22]~q ),
	.datac(\my_reg[8][22]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux9~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~12 .lut_mask = 16'hEE50;
defparam \Mux9~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N8
cycloneive_lcell_comb \Mux9~13 (
// Equation(s):
// \Mux9~13_combout  = (dcifimemload_21 & ((\Mux9~12_combout  & ((\my_reg[11][22]~q ))) # (!\Mux9~12_combout  & (\my_reg[9][22]~q )))) # (!dcifimemload_21 & (((\Mux9~12_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][22]~q ),
	.datac(\my_reg[11][22]~q ),
	.datad(\Mux9~12_combout ),
	.cin(gnd),
	.combout(\Mux9~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~13 .lut_mask = 16'hF588;
defparam \Mux9~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N16
cycloneive_lcell_comb \Mux9~16 (
// Equation(s):
// \Mux9~16_combout  = (dcifimemload_23 & (dcifimemload_24)) # (!dcifimemload_23 & ((dcifimemload_24 & ((\Mux9~13_combout ))) # (!dcifimemload_24 & (\Mux9~15_combout ))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux9~15_combout ),
	.datad(\Mux9~13_combout ),
	.cin(gnd),
	.combout(\Mux9~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~16 .lut_mask = 16'hDC98;
defparam \Mux9~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N8
cycloneive_lcell_comb \Mux9~19 (
// Equation(s):
// \Mux9~19_combout  = (dcifimemload_23 & ((\Mux9~16_combout  & (\Mux9~18_combout )) # (!\Mux9~16_combout  & ((\Mux9~11_combout ))))) # (!dcifimemload_23 & (((\Mux9~16_combout ))))

	.dataa(\Mux9~18_combout ),
	.datab(dcifimemload_23),
	.datac(\Mux9~11_combout ),
	.datad(\Mux9~16_combout ),
	.cin(gnd),
	.combout(\Mux9~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~19 .lut_mask = 16'hBBC0;
defparam \Mux9~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N19
dffeas \my_reg[23][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][22] .is_wysiwyg = "true";
defparam \my_reg[23][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y41_N23
dffeas \my_reg[31][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][22] .is_wysiwyg = "true";
defparam \my_reg[31][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y40_N5
dffeas \my_reg[27][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][22] .is_wysiwyg = "true";
defparam \my_reg[27][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y41_N25
dffeas \my_reg[19][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][22] .is_wysiwyg = "true";
defparam \my_reg[19][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N24
cycloneive_lcell_comb \Mux9~7 (
// Equation(s):
// \Mux9~7_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[27][22]~q )) # (!dcifimemload_24 & ((\my_reg[19][22]~q )))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[27][22]~q ),
	.datac(\my_reg[19][22]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux9~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~7 .lut_mask = 16'hEE50;
defparam \Mux9~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N22
cycloneive_lcell_comb \Mux9~8 (
// Equation(s):
// \Mux9~8_combout  = (dcifimemload_23 & ((\Mux9~7_combout  & ((\my_reg[31][22]~q ))) # (!\Mux9~7_combout  & (\my_reg[23][22]~q )))) # (!dcifimemload_23 & (((\Mux9~7_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[23][22]~q ),
	.datac(\my_reg[31][22]~q ),
	.datad(\Mux9~7_combout ),
	.cin(gnd),
	.combout(\Mux9~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~8 .lut_mask = 16'hF588;
defparam \Mux9~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N23
dffeas \my_reg[21][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][22] .is_wysiwyg = "true";
defparam \my_reg[21][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N25
dffeas \my_reg[29][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][22] .is_wysiwyg = "true";
defparam \my_reg[29][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N25
dffeas \my_reg[17][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][22] .is_wysiwyg = "true";
defparam \my_reg[17][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N24
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[25][22]~q )) # (!dcifimemload_24 & ((\my_reg[17][22]~q )))))

	.dataa(\my_reg[25][22]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[17][22]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hEE30;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N24
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// \Mux9~1_combout  = (dcifimemload_23 & ((\Mux9~0_combout  & ((\my_reg[29][22]~q ))) # (!\Mux9~0_combout  & (\my_reg[21][22]~q )))) # (!dcifimemload_23 & (((\Mux9~0_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[21][22]~q ),
	.datac(\my_reg[29][22]~q ),
	.datad(\Mux9~0_combout ),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hF588;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N15
dffeas \my_reg[30][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][22] .is_wysiwyg = "true";
defparam \my_reg[30][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N7
dffeas \my_reg[18][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][22] .is_wysiwyg = "true";
defparam \my_reg[18][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N12
cycloneive_lcell_comb \Mux9~2 (
// Equation(s):
// \Mux9~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[22][22]~q )) # (!dcifimemload_23 & ((\my_reg[18][22]~q )))))

	.dataa(\my_reg[22][22]~q ),
	.datab(\my_reg[18][22]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux9~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~2 .lut_mask = 16'hFA0C;
defparam \Mux9~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N14
cycloneive_lcell_comb \Mux9~3 (
// Equation(s):
// \Mux9~3_combout  = (dcifimemload_24 & ((\Mux9~2_combout  & ((\my_reg[30][22]~q ))) # (!\Mux9~2_combout  & (\my_reg[26][22]~q )))) # (!dcifimemload_24 & (((\Mux9~2_combout ))))

	.dataa(\my_reg[26][22]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[30][22]~q ),
	.datad(\Mux9~2_combout ),
	.cin(gnd),
	.combout(\Mux9~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~3 .lut_mask = 16'hF388;
defparam \Mux9~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y30_N7
dffeas \my_reg[28][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][22] .is_wysiwyg = "true";
defparam \my_reg[28][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N21
dffeas \my_reg[16][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][22] .is_wysiwyg = "true";
defparam \my_reg[16][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y42_N31
dffeas \my_reg[20][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][22] .is_wysiwyg = "true";
defparam \my_reg[20][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N20
cycloneive_lcell_comb \Mux9~4 (
// Equation(s):
// \Mux9~4_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & ((\my_reg[20][22]~q ))) # (!dcifimemload_23 & (\my_reg[16][22]~q ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\my_reg[16][22]~q ),
	.datad(\my_reg[20][22]~q ),
	.cin(gnd),
	.combout(\Mux9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~4 .lut_mask = 16'hDC98;
defparam \Mux9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N6
cycloneive_lcell_comb \Mux9~5 (
// Equation(s):
// \Mux9~5_combout  = (dcifimemload_24 & ((\Mux9~4_combout  & ((\my_reg[28][22]~q ))) # (!\Mux9~4_combout  & (\my_reg[24][22]~q )))) # (!dcifimemload_24 & (((\Mux9~4_combout ))))

	.dataa(\my_reg[24][22]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[28][22]~q ),
	.datad(\Mux9~4_combout ),
	.cin(gnd),
	.combout(\Mux9~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~5 .lut_mask = 16'hF388;
defparam \Mux9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N28
cycloneive_lcell_comb \Mux9~6 (
// Equation(s):
// \Mux9~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux9~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\Mux9~5_combout ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux9~3_combout ),
	.datad(\Mux9~5_combout ),
	.cin(gnd),
	.combout(\Mux9~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~6 .lut_mask = 16'hB9A8;
defparam \Mux9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N10
cycloneive_lcell_comb \Mux9~9 (
// Equation(s):
// \Mux9~9_combout  = (dcifimemload_21 & ((\Mux9~6_combout  & (\Mux9~8_combout )) # (!\Mux9~6_combout  & ((\Mux9~1_combout ))))) # (!dcifimemload_21 & (((\Mux9~6_combout ))))

	.dataa(\Mux9~8_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux9~1_combout ),
	.datad(\Mux9~6_combout ),
	.cin(gnd),
	.combout(\Mux9~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~9 .lut_mask = 16'hBBC0;
defparam \Mux9~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N2
cycloneive_lcell_comb \Mux41~0 (
// Equation(s):
// \Mux41~0_combout  = (dcifimemload_17 & (((\my_reg[10][22]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\my_reg[8][22]~q  & ((!dcifimemload_16))))

	.dataa(\my_reg[8][22]~q ),
	.datab(\my_reg[10][22]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux41~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~0 .lut_mask = 16'hF0CA;
defparam \Mux41~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N30
cycloneive_lcell_comb \Mux41~1 (
// Equation(s):
// \Mux41~1_combout  = (\Mux41~0_combout  & ((\my_reg[11][22]~q ) # ((!dcifimemload_16)))) # (!\Mux41~0_combout  & (((\my_reg[9][22]~q  & dcifimemload_16))))

	.dataa(\my_reg[11][22]~q ),
	.datab(\Mux41~0_combout ),
	.datac(\my_reg[9][22]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux41~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~1 .lut_mask = 16'hB8CC;
defparam \Mux41~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N26
cycloneive_lcell_comb \Mux41~5 (
// Equation(s):
// \Mux41~5_combout  = (\Mux41~4_combout ) # ((dcifimemload_17 & (\my_reg[2][22]~q  & !dcifimemload_16)))

	.dataa(\Mux41~4_combout ),
	.datab(dcifimemload_17),
	.datac(\my_reg[2][22]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux41~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~5 .lut_mask = 16'hAAEA;
defparam \Mux41~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N16
cycloneive_lcell_comb \Mux41~3 (
// Equation(s):
// \Mux41~3_combout  = (\Mux41~2_combout  & ((\my_reg[7][22]~q ) # ((!dcifimemload_17)))) # (!\Mux41~2_combout  & (((\my_reg[6][22]~q  & dcifimemload_17))))

	.dataa(\Mux41~2_combout ),
	.datab(\my_reg[7][22]~q ),
	.datac(\my_reg[6][22]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux41~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~3 .lut_mask = 16'hD8AA;
defparam \Mux41~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N4
cycloneive_lcell_comb \Mux41~6 (
// Equation(s):
// \Mux41~6_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & ((\Mux41~3_combout ))) # (!dcifimemload_18 & (\Mux41~5_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux41~5_combout ),
	.datad(\Mux41~3_combout ),
	.cin(gnd),
	.combout(\Mux41~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~6 .lut_mask = 16'hDC98;
defparam \Mux41~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N30
cycloneive_lcell_comb \Mux41~7 (
// Equation(s):
// \Mux41~7_combout  = (dcifimemload_16 & (((\my_reg[13][22]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[12][22]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[12][22]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[13][22]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux41~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~7 .lut_mask = 16'hCCE2;
defparam \Mux41~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N17
dffeas \my_reg[14][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][22] .is_wysiwyg = "true";
defparam \my_reg[14][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N16
cycloneive_lcell_comb \Mux41~8 (
// Equation(s):
// \Mux41~8_combout  = (\Mux41~7_combout  & ((\my_reg[15][22]~q ) # ((!dcifimemload_17)))) # (!\Mux41~7_combout  & (((\my_reg[14][22]~q  & dcifimemload_17))))

	.dataa(\Mux41~7_combout ),
	.datab(\my_reg[15][22]~q ),
	.datac(\my_reg[14][22]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux41~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~8 .lut_mask = 16'hD8AA;
defparam \Mux41~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N18
cycloneive_lcell_comb \Mux41~17 (
// Equation(s):
// \Mux41~17_combout  = (dcifimemload_18 & (((\my_reg[23][22]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[19][22]~q  & ((!dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[19][22]~q ),
	.datac(\my_reg[23][22]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux41~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~17 .lut_mask = 16'hAAE4;
defparam \Mux41~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N4
cycloneive_lcell_comb \Mux41~18 (
// Equation(s):
// \Mux41~18_combout  = (dcifimemload_19 & ((\Mux41~17_combout  & (\my_reg[31][22]~q )) # (!\Mux41~17_combout  & ((\my_reg[27][22]~q ))))) # (!dcifimemload_19 & (((\Mux41~17_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[31][22]~q ),
	.datac(\my_reg[27][22]~q ),
	.datad(\Mux41~17_combout ),
	.cin(gnd),
	.combout(\Mux41~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~18 .lut_mask = 16'hDDA0;
defparam \Mux41~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N6
cycloneive_lcell_comb \my_reg[25][22]~feeder (
// Equation(s):
// \my_reg[25][22]~feeder_combout  = \wdat~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat11),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[25][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][22]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[25][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N7
dffeas \my_reg[25][22] (
	.clk(CLK),
	.d(\my_reg[25][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][22] .is_wysiwyg = "true";
defparam \my_reg[25][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N10
cycloneive_lcell_comb \Mux41~10 (
// Equation(s):
// \Mux41~10_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[21][22]~q ))) # (!dcifimemload_18 & (\my_reg[17][22]~q ))))

	.dataa(\my_reg[17][22]~q ),
	.datab(\my_reg[21][22]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux41~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~10 .lut_mask = 16'hFC0A;
defparam \Mux41~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N28
cycloneive_lcell_comb \Mux41~11 (
// Equation(s):
// \Mux41~11_combout  = (dcifimemload_19 & ((\Mux41~10_combout  & ((\my_reg[29][22]~q ))) # (!\Mux41~10_combout  & (\my_reg[25][22]~q )))) # (!dcifimemload_19 & (((\Mux41~10_combout ))))

	.dataa(\my_reg[25][22]~q ),
	.datab(\my_reg[29][22]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux41~10_combout ),
	.cin(gnd),
	.combout(\Mux41~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~11 .lut_mask = 16'hCFA0;
defparam \Mux41~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y29_N25
dffeas \my_reg[24][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][22] .is_wysiwyg = "true";
defparam \my_reg[24][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N24
cycloneive_lcell_comb \Mux41~14 (
// Equation(s):
// \Mux41~14_combout  = (dcifimemload_19 & (((\my_reg[24][22]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[16][22]~q  & ((!dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[16][22]~q ),
	.datac(\my_reg[24][22]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux41~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~14 .lut_mask = 16'hAAE4;
defparam \Mux41~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N30
cycloneive_lcell_comb \Mux41~15 (
// Equation(s):
// \Mux41~15_combout  = (dcifimemload_18 & ((\Mux41~14_combout  & (\my_reg[28][22]~q )) # (!\Mux41~14_combout  & ((\my_reg[20][22]~q ))))) # (!dcifimemload_18 & (((\Mux41~14_combout ))))

	.dataa(\my_reg[28][22]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[20][22]~q ),
	.datad(\Mux41~14_combout ),
	.cin(gnd),
	.combout(\Mux41~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~15 .lut_mask = 16'hBBC0;
defparam \Mux41~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N11
dffeas \my_reg[22][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][22] .is_wysiwyg = "true";
defparam \my_reg[22][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N29
dffeas \my_reg[26][22] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][22] .is_wysiwyg = "true";
defparam \my_reg[26][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N28
cycloneive_lcell_comb \Mux41~12 (
// Equation(s):
// \Mux41~12_combout  = (dcifimemload_19 & (((\my_reg[26][22]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[18][22]~q  & ((!dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[18][22]~q ),
	.datac(\my_reg[26][22]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux41~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~12 .lut_mask = 16'hAAE4;
defparam \Mux41~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N10
cycloneive_lcell_comb \Mux41~13 (
// Equation(s):
// \Mux41~13_combout  = (dcifimemload_18 & ((\Mux41~12_combout  & (\my_reg[30][22]~q )) # (!\Mux41~12_combout  & ((\my_reg[22][22]~q ))))) # (!dcifimemload_18 & (((\Mux41~12_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[30][22]~q ),
	.datac(\my_reg[22][22]~q ),
	.datad(\Mux41~12_combout ),
	.cin(gnd),
	.combout(\Mux41~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~13 .lut_mask = 16'hDDA0;
defparam \Mux41~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N6
cycloneive_lcell_comb \Mux41~16 (
// Equation(s):
// \Mux41~16_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux41~13_combout ))) # (!dcifimemload_17 & (\Mux41~15_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux41~15_combout ),
	.datad(\Mux41~13_combout ),
	.cin(gnd),
	.combout(\Mux41~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~16 .lut_mask = 16'hDC98;
defparam \Mux41~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N31
dffeas \my_reg[2][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][21] .is_wysiwyg = "true";
defparam \my_reg[2][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N30
cycloneive_lcell_comb \Mux10~15 (
// Equation(s):
// \Mux10~15_combout  = (\Mux10~14_combout ) # ((!dcifimemload_21 & (\my_reg[2][21]~q  & dcifimemload_22)))

	.dataa(\Mux10~14_combout ),
	.datab(dcifimemload_21),
	.datac(\my_reg[2][21]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux10~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~15 .lut_mask = 16'hBAAA;
defparam \Mux10~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N9
dffeas \my_reg[6][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][21] .is_wysiwyg = "true";
defparam \my_reg[6][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N19
dffeas \my_reg[7][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][21] .is_wysiwyg = "true";
defparam \my_reg[7][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N30
cycloneive_lcell_comb \my_reg[4][21]~feeder (
// Equation(s):
// \my_reg[4][21]~feeder_combout  = \wdat~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat12),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[4][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[4][21]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[4][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N31
dffeas \my_reg[4][21] (
	.clk(CLK),
	.d(\my_reg[4][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][21] .is_wysiwyg = "true";
defparam \my_reg[4][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N28
cycloneive_lcell_comb \Mux10~12 (
// Equation(s):
// \Mux10~12_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\my_reg[5][21]~q )) # (!dcifimemload_21 & ((\my_reg[4][21]~q )))))

	.dataa(\my_reg[5][21]~q ),
	.datab(\my_reg[4][21]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux10~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~12 .lut_mask = 16'hFA0C;
defparam \Mux10~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N18
cycloneive_lcell_comb \Mux10~13 (
// Equation(s):
// \Mux10~13_combout  = (dcifimemload_22 & ((\Mux10~12_combout  & ((\my_reg[7][21]~q ))) # (!\Mux10~12_combout  & (\my_reg[6][21]~q )))) # (!dcifimemload_22 & (((\Mux10~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[6][21]~q ),
	.datac(\my_reg[7][21]~q ),
	.datad(\Mux10~12_combout ),
	.cin(gnd),
	.combout(\Mux10~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~13 .lut_mask = 16'hF588;
defparam \Mux10~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N4
cycloneive_lcell_comb \Mux10~16 (
// Equation(s):
// \Mux10~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & ((\Mux10~13_combout ))) # (!dcifimemload_23 & (\Mux10~15_combout ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux10~15_combout ),
	.datad(\Mux10~13_combout ),
	.cin(gnd),
	.combout(\Mux10~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~16 .lut_mask = 16'hDC98;
defparam \Mux10~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N31
dffeas \my_reg[15][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][21] .is_wysiwyg = "true";
defparam \my_reg[15][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y41_N21
dffeas \my_reg[14][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][21] .is_wysiwyg = "true";
defparam \my_reg[14][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N30
cycloneive_lcell_comb \Mux10~18 (
// Equation(s):
// \Mux10~18_combout  = (\Mux10~17_combout  & (((\my_reg[15][21]~q )) # (!dcifimemload_22))) # (!\Mux10~17_combout  & (dcifimemload_22 & ((\my_reg[14][21]~q ))))

	.dataa(\Mux10~17_combout ),
	.datab(dcifimemload_22),
	.datac(\my_reg[15][21]~q ),
	.datad(\my_reg[14][21]~q ),
	.cin(gnd),
	.combout(\Mux10~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~18 .lut_mask = 16'hE6A2;
defparam \Mux10~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y30_N25
dffeas \my_reg[9][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][21] .is_wysiwyg = "true";
defparam \my_reg[9][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y41_N11
dffeas \my_reg[11][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][21] .is_wysiwyg = "true";
defparam \my_reg[11][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N31
dffeas \my_reg[10][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][21] .is_wysiwyg = "true";
defparam \my_reg[10][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N14
cycloneive_lcell_comb \my_reg[8][21]~feeder (
// Equation(s):
// \my_reg[8][21]~feeder_combout  = \wdat~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat12),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[8][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[8][21]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[8][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N15
dffeas \my_reg[8][21] (
	.clk(CLK),
	.d(\my_reg[8][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][21] .is_wysiwyg = "true";
defparam \my_reg[8][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N16
cycloneive_lcell_comb \Mux10~10 (
// Equation(s):
// \Mux10~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][21]~q )) # (!dcifimemload_22 & ((\my_reg[8][21]~q )))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[10][21]~q ),
	.datac(\my_reg[8][21]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux10~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~10 .lut_mask = 16'hEE50;
defparam \Mux10~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N10
cycloneive_lcell_comb \Mux10~11 (
// Equation(s):
// \Mux10~11_combout  = (dcifimemload_21 & ((\Mux10~10_combout  & ((\my_reg[11][21]~q ))) # (!\Mux10~10_combout  & (\my_reg[9][21]~q )))) # (!dcifimemload_21 & (((\Mux10~10_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][21]~q ),
	.datac(\my_reg[11][21]~q ),
	.datad(\Mux10~10_combout ),
	.cin(gnd),
	.combout(\Mux10~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~11 .lut_mask = 16'hF588;
defparam \Mux10~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N14
cycloneive_lcell_comb \Mux10~19 (
// Equation(s):
// \Mux10~19_combout  = (dcifimemload_24 & ((\Mux10~16_combout  & (\Mux10~18_combout )) # (!\Mux10~16_combout  & ((\Mux10~11_combout ))))) # (!dcifimemload_24 & (\Mux10~16_combout ))

	.dataa(dcifimemload_24),
	.datab(\Mux10~16_combout ),
	.datac(\Mux10~18_combout ),
	.datad(\Mux10~11_combout ),
	.cin(gnd),
	.combout(\Mux10~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~19 .lut_mask = 16'hE6C4;
defparam \Mux10~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N7
dffeas \my_reg[27][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][21] .is_wysiwyg = "true";
defparam \my_reg[27][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N15
dffeas \my_reg[31][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][21] .is_wysiwyg = "true";
defparam \my_reg[31][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N1
dffeas \my_reg[19][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][21] .is_wysiwyg = "true";
defparam \my_reg[19][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N0
cycloneive_lcell_comb \Mux10~7 (
// Equation(s):
// \Mux10~7_combout  = (dcifimemload_23 & ((\my_reg[23][21]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[19][21]~q  & !dcifimemload_24))))

	.dataa(\my_reg[23][21]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[19][21]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux10~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~7 .lut_mask = 16'hCCB8;
defparam \Mux10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N14
cycloneive_lcell_comb \Mux10~8 (
// Equation(s):
// \Mux10~8_combout  = (dcifimemload_24 & ((\Mux10~7_combout  & ((\my_reg[31][21]~q ))) # (!\Mux10~7_combout  & (\my_reg[27][21]~q )))) # (!dcifimemload_24 & (((\Mux10~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[27][21]~q ),
	.datac(\my_reg[31][21]~q ),
	.datad(\Mux10~7_combout ),
	.cin(gnd),
	.combout(\Mux10~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~8 .lut_mask = 16'hF588;
defparam \Mux10~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y42_N31
dffeas \my_reg[25][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][21] .is_wysiwyg = "true";
defparam \my_reg[25][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N19
dffeas \my_reg[29][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][21] .is_wysiwyg = "true";
defparam \my_reg[29][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N13
dffeas \my_reg[21][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][21] .is_wysiwyg = "true";
defparam \my_reg[21][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N27
dffeas \my_reg[17][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][21] .is_wysiwyg = "true";
defparam \my_reg[17][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N26
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (dcifimemload_23 & ((\my_reg[21][21]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[17][21]~q  & !dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[21][21]~q ),
	.datac(\my_reg[17][21]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hAAD8;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N18
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// \Mux10~1_combout  = (dcifimemload_24 & ((\Mux10~0_combout  & ((\my_reg[29][21]~q ))) # (!\Mux10~0_combout  & (\my_reg[25][21]~q )))) # (!dcifimemload_24 & (((\Mux10~0_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[25][21]~q ),
	.datac(\my_reg[29][21]~q ),
	.datad(\Mux10~0_combout ),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hF588;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N20
cycloneive_lcell_comb \my_reg[30][21]~feeder (
// Equation(s):
// \my_reg[30][21]~feeder_combout  = \wdat~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat12),
	.cin(gnd),
	.combout(\my_reg[30][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[30][21]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[30][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y42_N21
dffeas \my_reg[30][21] (
	.clk(CLK),
	.d(\my_reg[30][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][21] .is_wysiwyg = "true";
defparam \my_reg[30][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N16
cycloneive_lcell_comb \my_reg[18][21]~feeder (
// Equation(s):
// \my_reg[18][21]~feeder_combout  = \wdat~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat12),
	.cin(gnd),
	.combout(\my_reg[18][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[18][21]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[18][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N17
dffeas \my_reg[18][21] (
	.clk(CLK),
	.d(\my_reg[18][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][21] .is_wysiwyg = "true";
defparam \my_reg[18][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y42_N15
dffeas \my_reg[26][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][21] .is_wysiwyg = "true";
defparam \my_reg[26][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N14
cycloneive_lcell_comb \Mux10~2 (
// Equation(s):
// \Mux10~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\my_reg[26][21]~q ))) # (!dcifimemload_24 & (\my_reg[18][21]~q ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[18][21]~q ),
	.datac(\my_reg[26][21]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~2 .lut_mask = 16'hFA44;
defparam \Mux10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N14
cycloneive_lcell_comb \Mux10~3 (
// Equation(s):
// \Mux10~3_combout  = (dcifimemload_23 & ((\Mux10~2_combout  & ((\my_reg[30][21]~q ))) # (!\Mux10~2_combout  & (\my_reg[22][21]~q )))) # (!dcifimemload_23 & (((\Mux10~2_combout ))))

	.dataa(\my_reg[22][21]~q ),
	.datab(\my_reg[30][21]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux10~2_combout ),
	.cin(gnd),
	.combout(\Mux10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~3 .lut_mask = 16'hCFA0;
defparam \Mux10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y29_N11
dffeas \my_reg[20][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][21] .is_wysiwyg = "true";
defparam \my_reg[20][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N23
dffeas \my_reg[28][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][21] .is_wysiwyg = "true";
defparam \my_reg[28][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N4
cycloneive_lcell_comb \my_reg[24][21]~feeder (
// Equation(s):
// \my_reg[24][21]~feeder_combout  = \wdat~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat12),
	.cin(gnd),
	.combout(\my_reg[24][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[24][21]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[24][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y29_N5
dffeas \my_reg[24][21] (
	.clk(CLK),
	.d(\my_reg[24][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][21] .is_wysiwyg = "true";
defparam \my_reg[24][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N10
cycloneive_lcell_comb \my_reg[16][21]~feeder (
// Equation(s):
// \my_reg[16][21]~feeder_combout  = \wdat~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat12),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[16][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[16][21]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[16][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N11
dffeas \my_reg[16][21] (
	.clk(CLK),
	.d(\my_reg[16][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][21] .is_wysiwyg = "true";
defparam \my_reg[16][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N28
cycloneive_lcell_comb \Mux10~4 (
// Equation(s):
// \Mux10~4_combout  = (dcifimemload_24 & ((\my_reg[24][21]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\my_reg[16][21]~q  & !dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[24][21]~q ),
	.datac(\my_reg[16][21]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~4 .lut_mask = 16'hAAD8;
defparam \Mux10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N22
cycloneive_lcell_comb \Mux10~5 (
// Equation(s):
// \Mux10~5_combout  = (dcifimemload_23 & ((\Mux10~4_combout  & ((\my_reg[28][21]~q ))) # (!\Mux10~4_combout  & (\my_reg[20][21]~q )))) # (!dcifimemload_23 & (((\Mux10~4_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[20][21]~q ),
	.datac(\my_reg[28][21]~q ),
	.datad(\Mux10~4_combout ),
	.cin(gnd),
	.combout(\Mux10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~5 .lut_mask = 16'hF588;
defparam \Mux10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N0
cycloneive_lcell_comb \Mux10~6 (
// Equation(s):
// \Mux10~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux10~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\Mux10~5_combout ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux10~3_combout ),
	.datad(\Mux10~5_combout ),
	.cin(gnd),
	.combout(\Mux10~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~6 .lut_mask = 16'hB9A8;
defparam \Mux10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N6
cycloneive_lcell_comb \Mux10~9 (
// Equation(s):
// \Mux10~9_combout  = (dcifimemload_21 & ((\Mux10~6_combout  & (\Mux10~8_combout )) # (!\Mux10~6_combout  & ((\Mux10~1_combout ))))) # (!dcifimemload_21 & (((\Mux10~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux10~8_combout ),
	.datac(\Mux10~1_combout ),
	.datad(\Mux10~6_combout ),
	.cin(gnd),
	.combout(\Mux10~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~9 .lut_mask = 16'hDDA0;
defparam \Mux10~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N13
dffeas \my_reg[3][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][21] .is_wysiwyg = "true";
defparam \my_reg[3][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N28
cycloneive_lcell_comb \Mux42~4 (
// Equation(s):
// \Mux42~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][21]~q ))) # (!dcifimemload_17 & (\my_reg[1][21]~q ))))

	.dataa(\my_reg[1][21]~q ),
	.datab(dcifimemload_17),
	.datac(\my_reg[3][21]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux42~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~4 .lut_mask = 16'hE200;
defparam \Mux42~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N22
cycloneive_lcell_comb \Mux42~5 (
// Equation(s):
// \Mux42~5_combout  = (\Mux42~4_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \my_reg[2][21]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\my_reg[2][21]~q ),
	.datad(\Mux42~4_combout ),
	.cin(gnd),
	.combout(\Mux42~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~5 .lut_mask = 16'hFF40;
defparam \Mux42~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N24
cycloneive_lcell_comb \Mux42~3 (
// Equation(s):
// \Mux42~3_combout  = (\Mux42~2_combout  & ((\my_reg[11][21]~q ) # ((!dcifimemload_16)))) # (!\Mux42~2_combout  & (((\my_reg[9][21]~q  & dcifimemload_16))))

	.dataa(\Mux42~2_combout ),
	.datab(\my_reg[11][21]~q ),
	.datac(\my_reg[9][21]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux42~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~3 .lut_mask = 16'hD8AA;
defparam \Mux42~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N12
cycloneive_lcell_comb \Mux42~6 (
// Equation(s):
// \Mux42~6_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & ((\Mux42~3_combout ))) # (!dcifimemload_19 & (\Mux42~5_combout ))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux42~5_combout ),
	.datad(\Mux42~3_combout ),
	.cin(gnd),
	.combout(\Mux42~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~6 .lut_mask = 16'hDC98;
defparam \Mux42~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N3
dffeas \my_reg[5][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][21] .is_wysiwyg = "true";
defparam \my_reg[5][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N2
cycloneive_lcell_comb \Mux42~0 (
// Equation(s):
// \Mux42~0_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][21]~q ))) # (!dcifimemload_16 & (\my_reg[4][21]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[4][21]~q ),
	.datac(\my_reg[5][21]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux42~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~0 .lut_mask = 16'hFA44;
defparam \Mux42~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N8
cycloneive_lcell_comb \Mux42~1 (
// Equation(s):
// \Mux42~1_combout  = (dcifimemload_17 & ((\Mux42~0_combout  & (\my_reg[7][21]~q )) # (!\Mux42~0_combout  & ((\my_reg[6][21]~q ))))) # (!dcifimemload_17 & (((\Mux42~0_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[7][21]~q ),
	.datac(\my_reg[6][21]~q ),
	.datad(\Mux42~0_combout ),
	.cin(gnd),
	.combout(\Mux42~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~1 .lut_mask = 16'hDDA0;
defparam \Mux42~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N25
dffeas \my_reg[13][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][21] .is_wysiwyg = "true";
defparam \my_reg[13][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N24
cycloneive_lcell_comb \Mux42~7 (
// Equation(s):
// \Mux42~7_combout  = (dcifimemload_16 & (((\my_reg[13][21]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[12][21]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[12][21]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[13][21]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux42~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~7 .lut_mask = 16'hCCE2;
defparam \Mux42~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N20
cycloneive_lcell_comb \Mux42~8 (
// Equation(s):
// \Mux42~8_combout  = (dcifimemload_17 & ((\Mux42~7_combout  & (\my_reg[15][21]~q )) # (!\Mux42~7_combout  & ((\my_reg[14][21]~q ))))) # (!dcifimemload_17 & (((\Mux42~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[15][21]~q ),
	.datac(\my_reg[14][21]~q ),
	.datad(\Mux42~7_combout ),
	.cin(gnd),
	.combout(\Mux42~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~8 .lut_mask = 16'hDDA0;
defparam \Mux42~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N30
cycloneive_lcell_comb \Mux42~10 (
// Equation(s):
// \Mux42~10_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[25][21]~q ))) # (!dcifimemload_19 & (\my_reg[17][21]~q ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[17][21]~q ),
	.datac(\my_reg[25][21]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux42~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~10 .lut_mask = 16'hFA44;
defparam \Mux42~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N12
cycloneive_lcell_comb \Mux42~11 (
// Equation(s):
// \Mux42~11_combout  = (dcifimemload_18 & ((\Mux42~10_combout  & (\my_reg[29][21]~q )) # (!\Mux42~10_combout  & ((\my_reg[21][21]~q ))))) # (!dcifimemload_18 & (((\Mux42~10_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[29][21]~q ),
	.datac(\my_reg[21][21]~q ),
	.datad(\Mux42~10_combout ),
	.cin(gnd),
	.combout(\Mux42~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~11 .lut_mask = 16'hDDA0;
defparam \Mux42~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N10
cycloneive_lcell_comb \Mux42~14 (
// Equation(s):
// \Mux42~14_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[20][21]~q ))) # (!dcifimemload_18 & (\my_reg[16][21]~q ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[16][21]~q ),
	.datac(\my_reg[20][21]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux42~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~14 .lut_mask = 16'hFA44;
defparam \Mux42~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N10
cycloneive_lcell_comb \Mux42~15 (
// Equation(s):
// \Mux42~15_combout  = (\Mux42~14_combout  & ((\my_reg[28][21]~q ) # ((!dcifimemload_19)))) # (!\Mux42~14_combout  & (((\my_reg[24][21]~q  & dcifimemload_19))))

	.dataa(\my_reg[28][21]~q ),
	.datab(\my_reg[24][21]~q ),
	.datac(\Mux42~14_combout ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux42~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~15 .lut_mask = 16'hACF0;
defparam \Mux42~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y42_N21
dffeas \my_reg[22][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][21] .is_wysiwyg = "true";
defparam \my_reg[22][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N20
cycloneive_lcell_comb \Mux42~12 (
// Equation(s):
// \Mux42~12_combout  = (dcifimemload_18 & (((\my_reg[22][21]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[18][21]~q  & ((!dcifimemload_19))))

	.dataa(\my_reg[18][21]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[22][21]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux42~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~12 .lut_mask = 16'hCCE2;
defparam \Mux42~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N14
cycloneive_lcell_comb \Mux42~13 (
// Equation(s):
// \Mux42~13_combout  = (dcifimemload_19 & ((\Mux42~12_combout  & (\my_reg[30][21]~q )) # (!\Mux42~12_combout  & ((\my_reg[26][21]~q ))))) # (!dcifimemload_19 & (((\Mux42~12_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[30][21]~q ),
	.datac(\my_reg[26][21]~q ),
	.datad(\Mux42~12_combout ),
	.cin(gnd),
	.combout(\Mux42~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~13 .lut_mask = 16'hDDA0;
defparam \Mux42~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N14
cycloneive_lcell_comb \Mux42~16 (
// Equation(s):
// \Mux42~16_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux42~13_combout ))) # (!dcifimemload_17 & (\Mux42~15_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux42~15_combout ),
	.datad(\Mux42~13_combout ),
	.cin(gnd),
	.combout(\Mux42~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~16 .lut_mask = 16'hDC98;
defparam \Mux42~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N9
dffeas \my_reg[23][21] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][21] .is_wysiwyg = "true";
defparam \my_reg[23][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N6
cycloneive_lcell_comb \Mux42~17 (
// Equation(s):
// \Mux42~17_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[27][21]~q ))) # (!dcifimemload_19 & (\my_reg[19][21]~q ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[19][21]~q ),
	.datac(\my_reg[27][21]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux42~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~17 .lut_mask = 16'hFA44;
defparam \Mux42~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N8
cycloneive_lcell_comb \Mux42~18 (
// Equation(s):
// \Mux42~18_combout  = (dcifimemload_18 & ((\Mux42~17_combout  & (\my_reg[31][21]~q )) # (!\Mux42~17_combout  & ((\my_reg[23][21]~q ))))) # (!dcifimemload_18 & (((\Mux42~17_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[31][21]~q ),
	.datac(\my_reg[23][21]~q ),
	.datad(\Mux42~17_combout ),
	.cin(gnd),
	.combout(\Mux42~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~18 .lut_mask = 16'hDDA0;
defparam \Mux42~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y40_N15
dffeas \my_reg[2][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][20] .is_wysiwyg = "true";
defparam \my_reg[2][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y40_N17
dffeas \my_reg[1][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][20] .is_wysiwyg = "true";
defparam \my_reg[1][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N16
cycloneive_lcell_comb \Mux11~14 (
// Equation(s):
// \Mux11~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\my_reg[3][20]~q )) # (!dcifimemload_22 & ((\my_reg[1][20]~q )))))

	.dataa(\my_reg[3][20]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[1][20]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux11~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~14 .lut_mask = 16'h88C0;
defparam \Mux11~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N14
cycloneive_lcell_comb \Mux11~15 (
// Equation(s):
// \Mux11~15_combout  = (\Mux11~14_combout ) # ((dcifimemload_22 & (!dcifimemload_21 & \my_reg[2][20]~q )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\my_reg[2][20]~q ),
	.datad(\Mux11~14_combout ),
	.cin(gnd),
	.combout(\Mux11~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~15 .lut_mask = 16'hFF20;
defparam \Mux11~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N4
cycloneive_lcell_comb \Mux11~16 (
// Equation(s):
// \Mux11~16_combout  = (dcifimemload_24 & ((\Mux11~13_combout ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\Mux11~15_combout  & !dcifimemload_23))))

	.dataa(\Mux11~13_combout ),
	.datab(dcifimemload_24),
	.datac(\Mux11~15_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux11~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~16 .lut_mask = 16'hCCB8;
defparam \Mux11~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N29
dffeas \my_reg[6][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][20] .is_wysiwyg = "true";
defparam \my_reg[6][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y42_N7
dffeas \my_reg[5][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][20] .is_wysiwyg = "true";
defparam \my_reg[5][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N17
dffeas \my_reg[4][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][20] .is_wysiwyg = "true";
defparam \my_reg[4][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N16
cycloneive_lcell_comb \Mux11~10 (
// Equation(s):
// \Mux11~10_combout  = (dcifimemload_21 & ((\my_reg[5][20]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[4][20]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[5][20]~q ),
	.datac(\my_reg[4][20]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux11~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~10 .lut_mask = 16'hAAD8;
defparam \Mux11~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N24
cycloneive_lcell_comb \Mux11~11 (
// Equation(s):
// \Mux11~11_combout  = (\Mux11~10_combout  & ((\my_reg[7][20]~q ) # ((!dcifimemload_22)))) # (!\Mux11~10_combout  & (((\my_reg[6][20]~q  & dcifimemload_22))))

	.dataa(\my_reg[7][20]~q ),
	.datab(\my_reg[6][20]~q ),
	.datac(\Mux11~10_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux11~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~11 .lut_mask = 16'hACF0;
defparam \Mux11~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N1
dffeas \my_reg[14][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][20] .is_wysiwyg = "true";
defparam \my_reg[14][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N3
dffeas \my_reg[15][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][20] .is_wysiwyg = "true";
defparam \my_reg[15][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N11
dffeas \my_reg[13][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][20] .is_wysiwyg = "true";
defparam \my_reg[13][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N11
dffeas \my_reg[12][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][20] .is_wysiwyg = "true";
defparam \my_reg[12][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N10
cycloneive_lcell_comb \Mux11~17 (
// Equation(s):
// \Mux11~17_combout  = (dcifimemload_21 & ((\my_reg[13][20]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][20]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[13][20]~q ),
	.datac(\my_reg[12][20]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux11~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~17 .lut_mask = 16'hAAD8;
defparam \Mux11~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N2
cycloneive_lcell_comb \Mux11~18 (
// Equation(s):
// \Mux11~18_combout  = (dcifimemload_22 & ((\Mux11~17_combout  & ((\my_reg[15][20]~q ))) # (!\Mux11~17_combout  & (\my_reg[14][20]~q )))) # (!dcifimemload_22 & (((\Mux11~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[14][20]~q ),
	.datac(\my_reg[15][20]~q ),
	.datad(\Mux11~17_combout ),
	.cin(gnd),
	.combout(\Mux11~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~18 .lut_mask = 16'hF588;
defparam \Mux11~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N22
cycloneive_lcell_comb \Mux11~19 (
// Equation(s):
// \Mux11~19_combout  = (dcifimemload_23 & ((\Mux11~16_combout  & ((\Mux11~18_combout ))) # (!\Mux11~16_combout  & (\Mux11~11_combout )))) # (!dcifimemload_23 & (\Mux11~16_combout ))

	.dataa(dcifimemload_23),
	.datab(\Mux11~16_combout ),
	.datac(\Mux11~11_combout ),
	.datad(\Mux11~18_combout ),
	.cin(gnd),
	.combout(\Mux11~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~19 .lut_mask = 16'hEC64;
defparam \Mux11~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N11
dffeas \my_reg[23][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][20] .is_wysiwyg = "true";
defparam \my_reg[23][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y41_N7
dffeas \my_reg[31][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][20] .is_wysiwyg = "true";
defparam \my_reg[31][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y40_N21
dffeas \my_reg[27][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][20] .is_wysiwyg = "true";
defparam \my_reg[27][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y41_N29
dffeas \my_reg[19][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][20] .is_wysiwyg = "true";
defparam \my_reg[19][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N28
cycloneive_lcell_comb \Mux11~7 (
// Equation(s):
// \Mux11~7_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[27][20]~q )) # (!dcifimemload_24 & ((\my_reg[19][20]~q )))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[27][20]~q ),
	.datac(\my_reg[19][20]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux11~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~7 .lut_mask = 16'hEE50;
defparam \Mux11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N6
cycloneive_lcell_comb \Mux11~8 (
// Equation(s):
// \Mux11~8_combout  = (dcifimemload_23 & ((\Mux11~7_combout  & ((\my_reg[31][20]~q ))) # (!\Mux11~7_combout  & (\my_reg[23][20]~q )))) # (!dcifimemload_23 & (((\Mux11~7_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[23][20]~q ),
	.datac(\my_reg[31][20]~q ),
	.datad(\Mux11~7_combout ),
	.cin(gnd),
	.combout(\Mux11~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~8 .lut_mask = 16'hF588;
defparam \Mux11~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N21
dffeas \my_reg[21][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][20] .is_wysiwyg = "true";
defparam \my_reg[21][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N7
dffeas \my_reg[17][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][20] .is_wysiwyg = "true";
defparam \my_reg[17][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N22
cycloneive_lcell_comb \my_reg[25][20]~feeder (
// Equation(s):
// \my_reg[25][20]~feeder_combout  = \wdat~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat13),
	.cin(gnd),
	.combout(\my_reg[25][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][20]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[25][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N23
dffeas \my_reg[25][20] (
	.clk(CLK),
	.d(\my_reg[25][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][20] .is_wysiwyg = "true";
defparam \my_reg[25][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N6
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (dcifimemload_24 & ((dcifimemload_23) # ((\my_reg[25][20]~q )))) # (!dcifimemload_24 & (!dcifimemload_23 & (\my_reg[17][20]~q )))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\my_reg[17][20]~q ),
	.datad(\my_reg[25][20]~q ),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hBA98;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N4
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// \Mux11~1_combout  = (dcifimemload_23 & ((\Mux11~0_combout  & (\my_reg[29][20]~q )) # (!\Mux11~0_combout  & ((\my_reg[21][20]~q ))))) # (!dcifimemload_23 & (((\Mux11~0_combout ))))

	.dataa(\my_reg[29][20]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[21][20]~q ),
	.datad(\Mux11~0_combout ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hBBC0;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N27
dffeas \my_reg[30][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][20] .is_wysiwyg = "true";
defparam \my_reg[30][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N19
dffeas \my_reg[18][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][20] .is_wysiwyg = "true";
defparam \my_reg[18][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N18
cycloneive_lcell_comb \Mux11~2 (
// Equation(s):
// \Mux11~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[22][20]~q )) # (!dcifimemload_23 & ((\my_reg[18][20]~q )))))

	.dataa(\my_reg[22][20]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[18][20]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~2 .lut_mask = 16'hEE30;
defparam \Mux11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N26
cycloneive_lcell_comb \Mux11~3 (
// Equation(s):
// \Mux11~3_combout  = (dcifimemload_24 & ((\Mux11~2_combout  & ((\my_reg[30][20]~q ))) # (!\Mux11~2_combout  & (\my_reg[26][20]~q )))) # (!dcifimemload_24 & (((\Mux11~2_combout ))))

	.dataa(\my_reg[26][20]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[30][20]~q ),
	.datad(\Mux11~2_combout ),
	.cin(gnd),
	.combout(\Mux11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~3 .lut_mask = 16'hF388;
defparam \Mux11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y32_N21
dffeas \my_reg[28][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][20] .is_wysiwyg = "true";
defparam \my_reg[28][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N3
dffeas \my_reg[20][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][20] .is_wysiwyg = "true";
defparam \my_reg[20][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N2
cycloneive_lcell_comb \Mux11~4 (
// Equation(s):
// \Mux11~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\my_reg[20][20]~q ))) # (!dcifimemload_23 & (\my_reg[16][20]~q ))))

	.dataa(\my_reg[16][20]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[20][20]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~4 .lut_mask = 16'hFC22;
defparam \Mux11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N16
cycloneive_lcell_comb \Mux11~5 (
// Equation(s):
// \Mux11~5_combout  = (dcifimemload_24 & ((\Mux11~4_combout  & ((\my_reg[28][20]~q ))) # (!\Mux11~4_combout  & (\my_reg[24][20]~q )))) # (!dcifimemload_24 & (((\Mux11~4_combout ))))

	.dataa(\my_reg[24][20]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[28][20]~q ),
	.datad(\Mux11~4_combout ),
	.cin(gnd),
	.combout(\Mux11~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~5 .lut_mask = 16'hF388;
defparam \Mux11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N24
cycloneive_lcell_comb \Mux11~6 (
// Equation(s):
// \Mux11~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux11~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\Mux11~5_combout ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux11~3_combout ),
	.datad(\Mux11~5_combout ),
	.cin(gnd),
	.combout(\Mux11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~6 .lut_mask = 16'hB9A8;
defparam \Mux11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N10
cycloneive_lcell_comb \Mux11~9 (
// Equation(s):
// \Mux11~9_combout  = (dcifimemload_21 & ((\Mux11~6_combout  & (\Mux11~8_combout )) # (!\Mux11~6_combout  & ((\Mux11~1_combout ))))) # (!dcifimemload_21 & (((\Mux11~6_combout ))))

	.dataa(\Mux11~8_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux11~1_combout ),
	.datad(\Mux11~6_combout ),
	.cin(gnd),
	.combout(\Mux11~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~9 .lut_mask = 16'hBBC0;
defparam \Mux11~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N5
dffeas \my_reg[8][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][20] .is_wysiwyg = "true";
defparam \my_reg[8][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N27
dffeas \my_reg[10][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][20] .is_wysiwyg = "true";
defparam \my_reg[10][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N26
cycloneive_lcell_comb \Mux43~0 (
// Equation(s):
// \Mux43~0_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[10][20]~q ))) # (!dcifimemload_17 & (\my_reg[8][20]~q ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[8][20]~q ),
	.datac(\my_reg[10][20]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux43~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~0 .lut_mask = 16'hFA44;
defparam \Mux43~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N23
dffeas \my_reg[11][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][20] .is_wysiwyg = "true";
defparam \my_reg[11][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N1
dffeas \my_reg[9][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][20] .is_wysiwyg = "true";
defparam \my_reg[9][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N0
cycloneive_lcell_comb \Mux43~1 (
// Equation(s):
// \Mux43~1_combout  = (\Mux43~0_combout  & ((\my_reg[11][20]~q ) # ((!dcifimemload_16)))) # (!\Mux43~0_combout  & (((\my_reg[9][20]~q  & dcifimemload_16))))

	.dataa(\Mux43~0_combout ),
	.datab(\my_reg[11][20]~q ),
	.datac(\my_reg[9][20]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux43~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~1 .lut_mask = 16'hD8AA;
defparam \Mux43~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N26
cycloneive_lcell_comb \my_reg[7][20]~feeder (
// Equation(s):
// \my_reg[7][20]~feeder_combout  = \wdat~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat13),
	.cin(gnd),
	.combout(\my_reg[7][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[7][20]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[7][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N27
dffeas \my_reg[7][20] (
	.clk(CLK),
	.d(\my_reg[7][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][20] .is_wysiwyg = "true";
defparam \my_reg[7][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N6
cycloneive_lcell_comb \Mux43~2 (
// Equation(s):
// \Mux43~2_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][20]~q ))) # (!dcifimemload_16 & (\my_reg[4][20]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[4][20]~q ),
	.datac(\my_reg[5][20]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux43~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~2 .lut_mask = 16'hFA44;
defparam \Mux43~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N28
cycloneive_lcell_comb \Mux43~3 (
// Equation(s):
// \Mux43~3_combout  = (dcifimemload_17 & ((\Mux43~2_combout  & (\my_reg[7][20]~q )) # (!\Mux43~2_combout  & ((\my_reg[6][20]~q ))))) # (!dcifimemload_17 & (((\Mux43~2_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[7][20]~q ),
	.datac(\my_reg[6][20]~q ),
	.datad(\Mux43~2_combout ),
	.cin(gnd),
	.combout(\Mux43~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~3 .lut_mask = 16'hDDA0;
defparam \Mux43~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N15
dffeas \my_reg[3][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][20] .is_wysiwyg = "true";
defparam \my_reg[3][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N14
cycloneive_lcell_comb \Mux43~4 (
// Equation(s):
// \Mux43~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][20]~q ))) # (!dcifimemload_17 & (\my_reg[1][20]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[1][20]~q ),
	.datac(\my_reg[3][20]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux43~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~4 .lut_mask = 16'hE400;
defparam \Mux43~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N0
cycloneive_lcell_comb \Mux43~5 (
// Equation(s):
// \Mux43~5_combout  = (\Mux43~4_combout ) # ((!dcifimemload_16 & (\my_reg[2][20]~q  & dcifimemload_17)))

	.dataa(dcifimemload_16),
	.datab(\my_reg[2][20]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux43~4_combout ),
	.cin(gnd),
	.combout(\Mux43~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~5 .lut_mask = 16'hFF40;
defparam \Mux43~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N26
cycloneive_lcell_comb \Mux43~6 (
// Equation(s):
// \Mux43~6_combout  = (dcifimemload_18 & ((dcifimemload_19) # ((\Mux43~3_combout )))) # (!dcifimemload_18 & (!dcifimemload_19 & ((\Mux43~5_combout ))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux43~3_combout ),
	.datad(\Mux43~5_combout ),
	.cin(gnd),
	.combout(\Mux43~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~6 .lut_mask = 16'hB9A8;
defparam \Mux43~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N10
cycloneive_lcell_comb \Mux43~7 (
// Equation(s):
// \Mux43~7_combout  = (dcifimemload_16 & (((\my_reg[13][20]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[12][20]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[12][20]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[13][20]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux43~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~7 .lut_mask = 16'hCCE2;
defparam \Mux43~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N0
cycloneive_lcell_comb \Mux43~8 (
// Equation(s):
// \Mux43~8_combout  = (dcifimemload_17 & ((\Mux43~7_combout  & (\my_reg[15][20]~q )) # (!\Mux43~7_combout  & ((\my_reg[14][20]~q ))))) # (!dcifimemload_17 & (((\Mux43~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[15][20]~q ),
	.datac(\my_reg[14][20]~q ),
	.datad(\Mux43~7_combout ),
	.cin(gnd),
	.combout(\Mux43~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~8 .lut_mask = 16'hDDA0;
defparam \Mux43~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N10
cycloneive_lcell_comb \Mux43~17 (
// Equation(s):
// \Mux43~17_combout  = (dcifimemload_18 & (((\my_reg[23][20]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[19][20]~q  & ((!dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[19][20]~q ),
	.datac(\my_reg[23][20]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux43~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~17 .lut_mask = 16'hAAE4;
defparam \Mux43~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N20
cycloneive_lcell_comb \Mux43~18 (
// Equation(s):
// \Mux43~18_combout  = (dcifimemload_19 & ((\Mux43~17_combout  & (\my_reg[31][20]~q )) # (!\Mux43~17_combout  & ((\my_reg[27][20]~q ))))) # (!dcifimemload_19 & (((\Mux43~17_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[31][20]~q ),
	.datac(\my_reg[27][20]~q ),
	.datad(\Mux43~17_combout ),
	.cin(gnd),
	.combout(\Mux43~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~18 .lut_mask = 16'hDDA0;
defparam \Mux43~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N20
cycloneive_lcell_comb \Mux43~10 (
// Equation(s):
// \Mux43~10_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[21][20]~q ))) # (!dcifimemload_18 & (\my_reg[17][20]~q ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[17][20]~q ),
	.datac(\my_reg[21][20]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux43~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~10 .lut_mask = 16'hFA44;
defparam \Mux43~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N6
cycloneive_lcell_comb \my_reg[29][20]~feeder (
// Equation(s):
// \my_reg[29][20]~feeder_combout  = \wdat~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat13),
	.cin(gnd),
	.combout(\my_reg[29][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[29][20]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[29][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N7
dffeas \my_reg[29][20] (
	.clk(CLK),
	.d(\my_reg[29][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][20] .is_wysiwyg = "true";
defparam \my_reg[29][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N14
cycloneive_lcell_comb \Mux43~11 (
// Equation(s):
// \Mux43~11_combout  = (dcifimemload_19 & ((\Mux43~10_combout  & ((\my_reg[29][20]~q ))) # (!\Mux43~10_combout  & (\my_reg[25][20]~q )))) # (!dcifimemload_19 & (((\Mux43~10_combout ))))

	.dataa(\my_reg[25][20]~q ),
	.datab(dcifimemload_19),
	.datac(\Mux43~10_combout ),
	.datad(\my_reg[29][20]~q ),
	.cin(gnd),
	.combout(\Mux43~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~11 .lut_mask = 16'hF838;
defparam \Mux43~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N23
dffeas \my_reg[16][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][20] .is_wysiwyg = "true";
defparam \my_reg[16][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N9
dffeas \my_reg[24][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][20] .is_wysiwyg = "true";
defparam \my_reg[24][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N8
cycloneive_lcell_comb \Mux43~14 (
// Equation(s):
// \Mux43~14_combout  = (dcifimemload_19 & (((\my_reg[24][20]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[16][20]~q  & ((!dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[16][20]~q ),
	.datac(\my_reg[24][20]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux43~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~14 .lut_mask = 16'hAAE4;
defparam \Mux43~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N26
cycloneive_lcell_comb \Mux43~15 (
// Equation(s):
// \Mux43~15_combout  = (\Mux43~14_combout  & ((\my_reg[28][20]~q ) # ((!dcifimemload_18)))) # (!\Mux43~14_combout  & (((\my_reg[20][20]~q  & dcifimemload_18))))

	.dataa(\my_reg[28][20]~q ),
	.datab(\Mux43~14_combout ),
	.datac(\my_reg[20][20]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux43~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~15 .lut_mask = 16'hB8CC;
defparam \Mux43~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N8
cycloneive_lcell_comb \my_reg[22][20]~feeder (
// Equation(s):
// \my_reg[22][20]~feeder_combout  = \wdat~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat13),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[22][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[22][20]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[22][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N9
dffeas \my_reg[22][20] (
	.clk(CLK),
	.d(\my_reg[22][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][20] .is_wysiwyg = "true";
defparam \my_reg[22][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N17
dffeas \my_reg[26][20] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][20] .is_wysiwyg = "true";
defparam \my_reg[26][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N16
cycloneive_lcell_comb \Mux43~12 (
// Equation(s):
// \Mux43~12_combout  = (dcifimemload_19 & (((\my_reg[26][20]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[18][20]~q  & ((!dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[18][20]~q ),
	.datac(\my_reg[26][20]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux43~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~12 .lut_mask = 16'hAAE4;
defparam \Mux43~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N24
cycloneive_lcell_comb \Mux43~13 (
// Equation(s):
// \Mux43~13_combout  = (dcifimemload_18 & ((\Mux43~12_combout  & (\my_reg[30][20]~q )) # (!\Mux43~12_combout  & ((\my_reg[22][20]~q ))))) # (!dcifimemload_18 & (((\Mux43~12_combout ))))

	.dataa(\my_reg[30][20]~q ),
	.datab(\my_reg[22][20]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux43~12_combout ),
	.cin(gnd),
	.combout(\Mux43~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~13 .lut_mask = 16'hAFC0;
defparam \Mux43~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N18
cycloneive_lcell_comb \Mux43~16 (
// Equation(s):
// \Mux43~16_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux43~13_combout ))) # (!dcifimemload_17 & (\Mux43~15_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux43~15_combout ),
	.datad(\Mux43~13_combout ),
	.cin(gnd),
	.combout(\Mux43~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~16 .lut_mask = 16'hDC98;
defparam \Mux43~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N9
dffeas \my_reg[19][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][19] .is_wysiwyg = "true";
defparam \my_reg[19][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N8
cycloneive_lcell_comb \Mux12~7 (
// Equation(s):
// \Mux12~7_combout  = (dcifimemload_23 & ((\my_reg[23][19]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[19][19]~q  & !dcifimemload_24))))

	.dataa(\my_reg[23][19]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[19][19]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux12~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~7 .lut_mask = 16'hCCB8;
defparam \Mux12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N19
dffeas \my_reg[31][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][19] .is_wysiwyg = "true";
defparam \my_reg[31][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N18
cycloneive_lcell_comb \Mux12~8 (
// Equation(s):
// \Mux12~8_combout  = (\Mux12~7_combout  & (((\my_reg[31][19]~q ) # (!dcifimemload_24)))) # (!\Mux12~7_combout  & (\my_reg[27][19]~q  & ((dcifimemload_24))))

	.dataa(\my_reg[27][19]~q ),
	.datab(\Mux12~7_combout ),
	.datac(\my_reg[31][19]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux12~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~8 .lut_mask = 16'hE2CC;
defparam \Mux12~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y30_N9
dffeas \my_reg[16][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][19] .is_wysiwyg = "true";
defparam \my_reg[16][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N8
cycloneive_lcell_comb \Mux12~4 (
// Equation(s):
// \Mux12~4_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[24][19]~q )) # (!dcifimemload_24 & ((\my_reg[16][19]~q )))))

	.dataa(\my_reg[24][19]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[16][19]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~4 .lut_mask = 16'hEE30;
defparam \Mux12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y30_N15
dffeas \my_reg[28][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][19] .is_wysiwyg = "true";
defparam \my_reg[28][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N14
cycloneive_lcell_comb \Mux12~5 (
// Equation(s):
// \Mux12~5_combout  = (\Mux12~4_combout  & (((\my_reg[28][19]~q ) # (!dcifimemload_23)))) # (!\Mux12~4_combout  & (\my_reg[20][19]~q  & ((dcifimemload_23))))

	.dataa(\my_reg[20][19]~q ),
	.datab(\Mux12~4_combout ),
	.datac(\my_reg[28][19]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux12~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~5 .lut_mask = 16'hE2CC;
defparam \Mux12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y42_N13
dffeas \my_reg[22][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][19] .is_wysiwyg = "true";
defparam \my_reg[22][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y42_N7
dffeas \my_reg[30][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][19] .is_wysiwyg = "true";
defparam \my_reg[30][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y42_N19
dffeas \my_reg[26][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][19] .is_wysiwyg = "true";
defparam \my_reg[26][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N12
cycloneive_lcell_comb \my_reg[18][19]~feeder (
// Equation(s):
// \my_reg[18][19]~feeder_combout  = \wdat~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat14),
	.cin(gnd),
	.combout(\my_reg[18][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[18][19]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[18][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N13
dffeas \my_reg[18][19] (
	.clk(CLK),
	.d(\my_reg[18][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][19] .is_wysiwyg = "true";
defparam \my_reg[18][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N22
cycloneive_lcell_comb \Mux12~2 (
// Equation(s):
// \Mux12~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[26][19]~q )) # (!dcifimemload_24 & ((\my_reg[18][19]~q )))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[26][19]~q ),
	.datac(\my_reg[18][19]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux12~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~2 .lut_mask = 16'hEE50;
defparam \Mux12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N6
cycloneive_lcell_comb \Mux12~3 (
// Equation(s):
// \Mux12~3_combout  = (dcifimemload_23 & ((\Mux12~2_combout  & ((\my_reg[30][19]~q ))) # (!\Mux12~2_combout  & (\my_reg[22][19]~q )))) # (!dcifimemload_23 & (((\Mux12~2_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[22][19]~q ),
	.datac(\my_reg[30][19]~q ),
	.datad(\Mux12~2_combout ),
	.cin(gnd),
	.combout(\Mux12~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~3 .lut_mask = 16'hF588;
defparam \Mux12~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N4
cycloneive_lcell_comb \Mux12~6 (
// Equation(s):
// \Mux12~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux12~3_combout ))) # (!dcifimemload_22 & (\Mux12~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux12~5_combout ),
	.datad(\Mux12~3_combout ),
	.cin(gnd),
	.combout(\Mux12~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~6 .lut_mask = 16'hDC98;
defparam \Mux12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N8
cycloneive_lcell_comb \my_reg[25][19]~feeder (
// Equation(s):
// \my_reg[25][19]~feeder_combout  = \wdat~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat14),
	.cin(gnd),
	.combout(\my_reg[25][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][19]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[25][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y42_N9
dffeas \my_reg[25][19] (
	.clk(CLK),
	.d(\my_reg[25][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][19] .is_wysiwyg = "true";
defparam \my_reg[25][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N3
dffeas \my_reg[29][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][19] .is_wysiwyg = "true";
defparam \my_reg[29][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N24
cycloneive_lcell_comb \my_reg[17][19]~feeder (
// Equation(s):
// \my_reg[17][19]~feeder_combout  = \wdat~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat14),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[17][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[17][19]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[17][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N25
dffeas \my_reg[17][19] (
	.clk(CLK),
	.d(\my_reg[17][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][19] .is_wysiwyg = "true";
defparam \my_reg[17][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N30
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (dcifimemload_23 & ((\my_reg[21][19]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[17][19]~q  & !dcifimemload_24))))

	.dataa(\my_reg[21][19]~q ),
	.datab(\my_reg[17][19]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hF0AC;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N2
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// \Mux12~1_combout  = (dcifimemload_24 & ((\Mux12~0_combout  & ((\my_reg[29][19]~q ))) # (!\Mux12~0_combout  & (\my_reg[25][19]~q )))) # (!dcifimemload_24 & (((\Mux12~0_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[25][19]~q ),
	.datac(\my_reg[29][19]~q ),
	.datad(\Mux12~0_combout ),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hF588;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N30
cycloneive_lcell_comb \Mux12~9 (
// Equation(s):
// \Mux12~9_combout  = (dcifimemload_21 & ((\Mux12~6_combout  & (\Mux12~8_combout )) # (!\Mux12~6_combout  & ((\Mux12~1_combout ))))) # (!dcifimemload_21 & (((\Mux12~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux12~8_combout ),
	.datac(\Mux12~6_combout ),
	.datad(\Mux12~1_combout ),
	.cin(gnd),
	.combout(\Mux12~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~9 .lut_mask = 16'hDAD0;
defparam \Mux12~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N11
dffeas \my_reg[15][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][19] .is_wysiwyg = "true";
defparam \my_reg[15][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N29
dffeas \my_reg[13][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][19] .is_wysiwyg = "true";
defparam \my_reg[13][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N27
dffeas \my_reg[12][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][19] .is_wysiwyg = "true";
defparam \my_reg[12][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N26
cycloneive_lcell_comb \Mux12~17 (
// Equation(s):
// \Mux12~17_combout  = (dcifimemload_21 & ((\my_reg[13][19]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][19]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[13][19]~q ),
	.datac(\my_reg[12][19]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux12~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~17 .lut_mask = 16'hAAD8;
defparam \Mux12~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N22
cycloneive_lcell_comb \Mux12~18 (
// Equation(s):
// \Mux12~18_combout  = (dcifimemload_22 & ((\Mux12~17_combout  & ((\my_reg[15][19]~q ))) # (!\Mux12~17_combout  & (\my_reg[14][19]~q )))) # (!dcifimemload_22 & (((\Mux12~17_combout ))))

	.dataa(\my_reg[14][19]~q ),
	.datab(\my_reg[15][19]~q ),
	.datac(dcifimemload_22),
	.datad(\Mux12~17_combout ),
	.cin(gnd),
	.combout(\Mux12~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~18 .lut_mask = 16'hCFA0;
defparam \Mux12~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y30_N9
dffeas \my_reg[9][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][19] .is_wysiwyg = "true";
defparam \my_reg[9][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N1
dffeas \my_reg[11][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][19] .is_wysiwyg = "true";
defparam \my_reg[11][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N1
dffeas \my_reg[8][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][19] .is_wysiwyg = "true";
defparam \my_reg[8][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N0
cycloneive_lcell_comb \Mux12~10 (
// Equation(s):
// \Mux12~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][19]~q )) # (!dcifimemload_22 & ((\my_reg[8][19]~q )))))

	.dataa(\my_reg[10][19]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[8][19]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux12~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~10 .lut_mask = 16'hEE30;
defparam \Mux12~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N0
cycloneive_lcell_comb \Mux12~11 (
// Equation(s):
// \Mux12~11_combout  = (dcifimemload_21 & ((\Mux12~10_combout  & ((\my_reg[11][19]~q ))) # (!\Mux12~10_combout  & (\my_reg[9][19]~q )))) # (!dcifimemload_21 & (((\Mux12~10_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][19]~q ),
	.datac(\my_reg[11][19]~q ),
	.datad(\Mux12~10_combout ),
	.cin(gnd),
	.combout(\Mux12~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~11 .lut_mask = 16'hF588;
defparam \Mux12~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y43_N9
dffeas \my_reg[7][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][19] .is_wysiwyg = "true";
defparam \my_reg[7][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y42_N31
dffeas \my_reg[5][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][19] .is_wysiwyg = "true";
defparam \my_reg[5][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N1
dffeas \my_reg[4][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][19] .is_wysiwyg = "true";
defparam \my_reg[4][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N0
cycloneive_lcell_comb \Mux12~12 (
// Equation(s):
// \Mux12~12_combout  = (dcifimemload_21 & ((\my_reg[5][19]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[4][19]~q  & !dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[5][19]~q ),
	.datac(\my_reg[4][19]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux12~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~12 .lut_mask = 16'hAAD8;
defparam \Mux12~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N8
cycloneive_lcell_comb \Mux12~13 (
// Equation(s):
// \Mux12~13_combout  = (dcifimemload_22 & ((\Mux12~12_combout  & ((\my_reg[7][19]~q ))) # (!\Mux12~12_combout  & (\my_reg[6][19]~q )))) # (!dcifimemload_22 & (((\Mux12~12_combout ))))

	.dataa(\my_reg[6][19]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[7][19]~q ),
	.datad(\Mux12~12_combout ),
	.cin(gnd),
	.combout(\Mux12~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~13 .lut_mask = 16'hF388;
defparam \Mux12~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y43_N3
dffeas \my_reg[2][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][19] .is_wysiwyg = "true";
defparam \my_reg[2][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N11
dffeas \my_reg[1][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][19] .is_wysiwyg = "true";
defparam \my_reg[1][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N10
cycloneive_lcell_comb \Mux12~14 (
// Equation(s):
// \Mux12~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\my_reg[3][19]~q )) # (!dcifimemload_22 & ((\my_reg[1][19]~q )))))

	.dataa(\my_reg[3][19]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[1][19]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux12~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~14 .lut_mask = 16'h88C0;
defparam \Mux12~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N2
cycloneive_lcell_comb \Mux12~15 (
// Equation(s):
// \Mux12~15_combout  = (\Mux12~14_combout ) # ((!dcifimemload_21 & (dcifimemload_22 & \my_reg[2][19]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\my_reg[2][19]~q ),
	.datad(\Mux12~14_combout ),
	.cin(gnd),
	.combout(\Mux12~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~15 .lut_mask = 16'hFF40;
defparam \Mux12~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N12
cycloneive_lcell_comb \Mux12~16 (
// Equation(s):
// \Mux12~16_combout  = (dcifimemload_23 & ((dcifimemload_24) # ((\Mux12~13_combout )))) # (!dcifimemload_23 & (!dcifimemload_24 & ((\Mux12~15_combout ))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux12~13_combout ),
	.datad(\Mux12~15_combout ),
	.cin(gnd),
	.combout(\Mux12~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~16 .lut_mask = 16'hB9A8;
defparam \Mux12~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N6
cycloneive_lcell_comb \Mux12~19 (
// Equation(s):
// \Mux12~19_combout  = (dcifimemload_24 & ((\Mux12~16_combout  & (\Mux12~18_combout )) # (!\Mux12~16_combout  & ((\Mux12~11_combout ))))) # (!dcifimemload_24 & (((\Mux12~16_combout ))))

	.dataa(dcifimemload_24),
	.datab(\Mux12~18_combout ),
	.datac(\Mux12~11_combout ),
	.datad(\Mux12~16_combout ),
	.cin(gnd),
	.combout(\Mux12~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~19 .lut_mask = 16'hDDA0;
defparam \Mux12~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y30_N19
dffeas \my_reg[10][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][19] .is_wysiwyg = "true";
defparam \my_reg[10][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N18
cycloneive_lcell_comb \Mux44~2 (
// Equation(s):
// \Mux44~2_combout  = (dcifimemload_17 & (((\my_reg[10][19]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\my_reg[8][19]~q  & ((!dcifimemload_16))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[8][19]~q ),
	.datac(\my_reg[10][19]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux44~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~2 .lut_mask = 16'hAAE4;
defparam \Mux44~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N8
cycloneive_lcell_comb \Mux44~3 (
// Equation(s):
// \Mux44~3_combout  = (dcifimemload_16 & ((\Mux44~2_combout  & (\my_reg[11][19]~q )) # (!\Mux44~2_combout  & ((\my_reg[9][19]~q ))))) # (!dcifimemload_16 & (((\Mux44~2_combout ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[11][19]~q ),
	.datac(\my_reg[9][19]~q ),
	.datad(\Mux44~2_combout ),
	.cin(gnd),
	.combout(\Mux44~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~3 .lut_mask = 16'hDDA0;
defparam \Mux44~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N12
cycloneive_lcell_comb \my_reg[3][19]~feeder (
// Equation(s):
// \my_reg[3][19]~feeder_combout  = \wdat~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat14),
	.cin(gnd),
	.combout(\my_reg[3][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[3][19]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[3][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N13
dffeas \my_reg[3][19] (
	.clk(CLK),
	.d(\my_reg[3][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][19] .is_wysiwyg = "true";
defparam \my_reg[3][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N24
cycloneive_lcell_comb \Mux44~4 (
// Equation(s):
// \Mux44~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][19]~q ))) # (!dcifimemload_17 & (\my_reg[1][19]~q ))))

	.dataa(\my_reg[1][19]~q ),
	.datab(\my_reg[3][19]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux44~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~4 .lut_mask = 16'hCA00;
defparam \Mux44~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N28
cycloneive_lcell_comb \Mux44~5 (
// Equation(s):
// \Mux44~5_combout  = (\Mux44~4_combout ) # ((!dcifimemload_16 & (\my_reg[2][19]~q  & dcifimemload_17)))

	.dataa(dcifimemload_16),
	.datab(\my_reg[2][19]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux44~4_combout ),
	.cin(gnd),
	.combout(\Mux44~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~5 .lut_mask = 16'hFF40;
defparam \Mux44~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N10
cycloneive_lcell_comb \Mux44~6 (
// Equation(s):
// \Mux44~6_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\Mux44~3_combout )))) # (!dcifimemload_19 & (!dcifimemload_18 & ((\Mux44~5_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux44~3_combout ),
	.datad(\Mux44~5_combout ),
	.cin(gnd),
	.combout(\Mux44~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~6 .lut_mask = 16'hB9A8;
defparam \Mux44~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N12
cycloneive_lcell_comb \my_reg[14][19]~feeder (
// Equation(s):
// \my_reg[14][19]~feeder_combout  = \wdat~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat14),
	.cin(gnd),
	.combout(\my_reg[14][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[14][19]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[14][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N13
dffeas \my_reg[14][19] (
	.clk(CLK),
	.d(\my_reg[14][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][19] .is_wysiwyg = "true";
defparam \my_reg[14][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N28
cycloneive_lcell_comb \Mux44~7 (
// Equation(s):
// \Mux44~7_combout  = (dcifimemload_16 & (((\my_reg[13][19]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[12][19]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[12][19]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[13][19]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux44~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~7 .lut_mask = 16'hCCE2;
defparam \Mux44~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N12
cycloneive_lcell_comb \Mux44~8 (
// Equation(s):
// \Mux44~8_combout  = (dcifimemload_17 & ((\Mux44~7_combout  & ((\my_reg[15][19]~q ))) # (!\Mux44~7_combout  & (\my_reg[14][19]~q )))) # (!dcifimemload_17 & (((\Mux44~7_combout ))))

	.dataa(\my_reg[14][19]~q ),
	.datab(\my_reg[15][19]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux44~7_combout ),
	.cin(gnd),
	.combout(\Mux44~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~8 .lut_mask = 16'hCFA0;
defparam \Mux44~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N30
cycloneive_lcell_comb \Mux44~0 (
// Equation(s):
// \Mux44~0_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][19]~q ))) # (!dcifimemload_16 & (\my_reg[4][19]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[4][19]~q ),
	.datac(\my_reg[5][19]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux44~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~0 .lut_mask = 16'hFA44;
defparam \Mux44~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N21
dffeas \my_reg[6][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][19] .is_wysiwyg = "true";
defparam \my_reg[6][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N20
cycloneive_lcell_comb \Mux44~1 (
// Equation(s):
// \Mux44~1_combout  = (\Mux44~0_combout  & ((\my_reg[7][19]~q ) # ((!dcifimemload_17)))) # (!\Mux44~0_combout  & (((\my_reg[6][19]~q  & dcifimemload_17))))

	.dataa(\Mux44~0_combout ),
	.datab(\my_reg[7][19]~q ),
	.datac(\my_reg[6][19]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux44~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~1 .lut_mask = 16'hD8AA;
defparam \Mux44~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N21
dffeas \my_reg[21][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][19] .is_wysiwyg = "true";
defparam \my_reg[21][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N16
cycloneive_lcell_comb \Mux44~10 (
// Equation(s):
// \Mux44~10_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[25][19]~q ))) # (!dcifimemload_19 & (\my_reg[17][19]~q ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[17][19]~q ),
	.datac(\my_reg[25][19]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux44~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~10 .lut_mask = 16'hFA44;
defparam \Mux44~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N20
cycloneive_lcell_comb \Mux44~11 (
// Equation(s):
// \Mux44~11_combout  = (dcifimemload_18 & ((\Mux44~10_combout  & (\my_reg[29][19]~q )) # (!\Mux44~10_combout  & ((\my_reg[21][19]~q ))))) # (!dcifimemload_18 & (((\Mux44~10_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[29][19]~q ),
	.datac(\my_reg[21][19]~q ),
	.datad(\Mux44~10_combout ),
	.cin(gnd),
	.combout(\Mux44~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~11 .lut_mask = 16'hDDA0;
defparam \Mux44~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N0
cycloneive_lcell_comb \Mux44~17 (
// Equation(s):
// \Mux44~17_combout  = (dcifimemload_19 & ((\my_reg[27][19]~q ) # ((dcifimemload_18)))) # (!dcifimemload_19 & (((\my_reg[19][19]~q  & !dcifimemload_18))))

	.dataa(\my_reg[27][19]~q ),
	.datab(\my_reg[19][19]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux44~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~17 .lut_mask = 16'hF0AC;
defparam \Mux44~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N10
cycloneive_lcell_comb \my_reg[23][19]~feeder (
// Equation(s):
// \my_reg[23][19]~feeder_combout  = \wdat~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat14),
	.cin(gnd),
	.combout(\my_reg[23][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[23][19]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[23][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N11
dffeas \my_reg[23][19] (
	.clk(CLK),
	.d(\my_reg[23][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][19] .is_wysiwyg = "true";
defparam \my_reg[23][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N22
cycloneive_lcell_comb \Mux44~18 (
// Equation(s):
// \Mux44~18_combout  = (\Mux44~17_combout  & ((\my_reg[31][19]~q ) # ((!dcifimemload_18)))) # (!\Mux44~17_combout  & (((\my_reg[23][19]~q  & dcifimemload_18))))

	.dataa(\my_reg[31][19]~q ),
	.datab(\Mux44~17_combout ),
	.datac(\my_reg[23][19]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux44~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~18 .lut_mask = 16'hB8CC;
defparam \Mux44~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y29_N15
dffeas \my_reg[24][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][19] .is_wysiwyg = "true";
defparam \my_reg[24][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N1
dffeas \my_reg[20][19] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][19] .is_wysiwyg = "true";
defparam \my_reg[20][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N0
cycloneive_lcell_comb \Mux44~14 (
// Equation(s):
// \Mux44~14_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[20][19]~q ))) # (!dcifimemload_18 & (\my_reg[16][19]~q ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[16][19]~q ),
	.datac(\my_reg[20][19]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux44~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~14 .lut_mask = 16'hFA44;
defparam \Mux44~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N14
cycloneive_lcell_comb \Mux44~15 (
// Equation(s):
// \Mux44~15_combout  = (dcifimemload_19 & ((\Mux44~14_combout  & (\my_reg[28][19]~q )) # (!\Mux44~14_combout  & ((\my_reg[24][19]~q ))))) # (!dcifimemload_19 & (((\Mux44~14_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[28][19]~q ),
	.datac(\my_reg[24][19]~q ),
	.datad(\Mux44~14_combout ),
	.cin(gnd),
	.combout(\Mux44~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~15 .lut_mask = 16'hDDA0;
defparam \Mux44~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N12
cycloneive_lcell_comb \Mux44~12 (
// Equation(s):
// \Mux44~12_combout  = (dcifimemload_18 & (((\my_reg[22][19]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[18][19]~q  & ((!dcifimemload_19))))

	.dataa(\my_reg[18][19]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[22][19]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux44~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~12 .lut_mask = 16'hCCE2;
defparam \Mux44~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N18
cycloneive_lcell_comb \Mux44~13 (
// Equation(s):
// \Mux44~13_combout  = (dcifimemload_19 & ((\Mux44~12_combout  & (\my_reg[30][19]~q )) # (!\Mux44~12_combout  & ((\my_reg[26][19]~q ))))) # (!dcifimemload_19 & (((\Mux44~12_combout ))))

	.dataa(\my_reg[30][19]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[26][19]~q ),
	.datad(\Mux44~12_combout ),
	.cin(gnd),
	.combout(\Mux44~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~13 .lut_mask = 16'hBBC0;
defparam \Mux44~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N2
cycloneive_lcell_comb \Mux44~16 (
// Equation(s):
// \Mux44~16_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux44~13_combout ))) # (!dcifimemload_17 & (\Mux44~15_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux44~15_combout ),
	.datad(\Mux44~13_combout ),
	.cin(gnd),
	.combout(\Mux44~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~16 .lut_mask = 16'hDC98;
defparam \Mux44~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N31
dffeas \my_reg[15][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][18] .is_wysiwyg = "true";
defparam \my_reg[15][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N23
dffeas \my_reg[14][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][18] .is_wysiwyg = "true";
defparam \my_reg[14][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N1
dffeas \my_reg[12][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][18] .is_wysiwyg = "true";
defparam \my_reg[12][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N0
cycloneive_lcell_comb \Mux13~17 (
// Equation(s):
// \Mux13~17_combout  = (dcifimemload_21 & ((\my_reg[13][18]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][18]~q  & !dcifimemload_22))))

	.dataa(\my_reg[13][18]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[12][18]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux13~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~17 .lut_mask = 16'hCCB8;
defparam \Mux13~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N22
cycloneive_lcell_comb \Mux13~18 (
// Equation(s):
// \Mux13~18_combout  = (dcifimemload_22 & ((\Mux13~17_combout  & (\my_reg[15][18]~q )) # (!\Mux13~17_combout  & ((\my_reg[14][18]~q ))))) # (!dcifimemload_22 & (((\Mux13~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[15][18]~q ),
	.datac(\my_reg[14][18]~q ),
	.datad(\Mux13~17_combout ),
	.cin(gnd),
	.combout(\Mux13~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~18 .lut_mask = 16'hDDA0;
defparam \Mux13~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N9
dffeas \my_reg[4][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][18] .is_wysiwyg = "true";
defparam \my_reg[4][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N8
cycloneive_lcell_comb \Mux13~10 (
// Equation(s):
// \Mux13~10_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\my_reg[5][18]~q )) # (!dcifimemload_21 & ((\my_reg[4][18]~q )))))

	.dataa(\my_reg[5][18]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[4][18]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux13~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~10 .lut_mask = 16'hEE30;
defparam \Mux13~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N23
dffeas \my_reg[7][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][18] .is_wysiwyg = "true";
defparam \my_reg[7][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N22
cycloneive_lcell_comb \Mux13~11 (
// Equation(s):
// \Mux13~11_combout  = (\Mux13~10_combout  & (((\my_reg[7][18]~q ) # (!dcifimemload_22)))) # (!\Mux13~10_combout  & (\my_reg[6][18]~q  & ((dcifimemload_22))))

	.dataa(\my_reg[6][18]~q ),
	.datab(\Mux13~10_combout ),
	.datac(\my_reg[7][18]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux13~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~11 .lut_mask = 16'hE2CC;
defparam \Mux13~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N21
dffeas \my_reg[2][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][18] .is_wysiwyg = "true";
defparam \my_reg[2][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N11
dffeas \my_reg[1][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][18] .is_wysiwyg = "true";
defparam \my_reg[1][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N10
cycloneive_lcell_comb \Mux13~14 (
// Equation(s):
// \Mux13~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\my_reg[3][18]~q )) # (!dcifimemload_22 & ((\my_reg[1][18]~q )))))

	.dataa(\my_reg[3][18]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[1][18]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux13~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~14 .lut_mask = 16'h88C0;
defparam \Mux13~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N20
cycloneive_lcell_comb \Mux13~15 (
// Equation(s):
// \Mux13~15_combout  = (\Mux13~14_combout ) # ((dcifimemload_22 & (!dcifimemload_21 & \my_reg[2][18]~q )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\my_reg[2][18]~q ),
	.datad(\Mux13~14_combout ),
	.cin(gnd),
	.combout(\Mux13~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~15 .lut_mask = 16'hFF20;
defparam \Mux13~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y30_N23
dffeas \my_reg[9][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][18] .is_wysiwyg = "true";
defparam \my_reg[9][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N5
dffeas \my_reg[11][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][18] .is_wysiwyg = "true";
defparam \my_reg[11][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N11
dffeas \my_reg[8][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][18] .is_wysiwyg = "true";
defparam \my_reg[8][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N10
cycloneive_lcell_comb \Mux13~12 (
// Equation(s):
// \Mux13~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][18]~q )) # (!dcifimemload_22 & ((\my_reg[8][18]~q )))))

	.dataa(\my_reg[10][18]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[8][18]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux13~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~12 .lut_mask = 16'hEE30;
defparam \Mux13~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N4
cycloneive_lcell_comb \Mux13~13 (
// Equation(s):
// \Mux13~13_combout  = (dcifimemload_21 & ((\Mux13~12_combout  & ((\my_reg[11][18]~q ))) # (!\Mux13~12_combout  & (\my_reg[9][18]~q )))) # (!dcifimemload_21 & (((\Mux13~12_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][18]~q ),
	.datac(\my_reg[11][18]~q ),
	.datad(\Mux13~12_combout ),
	.cin(gnd),
	.combout(\Mux13~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~13 .lut_mask = 16'hF588;
defparam \Mux13~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N6
cycloneive_lcell_comb \Mux13~16 (
// Equation(s):
// \Mux13~16_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\Mux13~13_combout ))) # (!dcifimemload_24 & (\Mux13~15_combout ))))

	.dataa(dcifimemload_23),
	.datab(\Mux13~15_combout ),
	.datac(dcifimemload_24),
	.datad(\Mux13~13_combout ),
	.cin(gnd),
	.combout(\Mux13~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~16 .lut_mask = 16'hF4A4;
defparam \Mux13~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N8
cycloneive_lcell_comb \Mux13~19 (
// Equation(s):
// \Mux13~19_combout  = (dcifimemload_23 & ((\Mux13~16_combout  & (\Mux13~18_combout )) # (!\Mux13~16_combout  & ((\Mux13~11_combout ))))) # (!dcifimemload_23 & (((\Mux13~16_combout ))))

	.dataa(dcifimemload_23),
	.datab(\Mux13~18_combout ),
	.datac(\Mux13~11_combout ),
	.datad(\Mux13~16_combout ),
	.cin(gnd),
	.combout(\Mux13~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~19 .lut_mask = 16'hDDA0;
defparam \Mux13~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N27
dffeas \my_reg[27][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][18] .is_wysiwyg = "true";
defparam \my_reg[27][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y41_N5
dffeas \my_reg[19][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][18] .is_wysiwyg = "true";
defparam \my_reg[19][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N4
cycloneive_lcell_comb \Mux13~7 (
// Equation(s):
// \Mux13~7_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[27][18]~q )) # (!dcifimemload_24 & ((\my_reg[19][18]~q )))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[27][18]~q ),
	.datac(\my_reg[19][18]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux13~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~7 .lut_mask = 16'hEE50;
defparam \Mux13~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N27
dffeas \my_reg[31][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][18] .is_wysiwyg = "true";
defparam \my_reg[31][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N26
cycloneive_lcell_comb \Mux13~8 (
// Equation(s):
// \Mux13~8_combout  = (\Mux13~7_combout  & (((\my_reg[31][18]~q ) # (!dcifimemload_23)))) # (!\Mux13~7_combout  & (\my_reg[23][18]~q  & ((dcifimemload_23))))

	.dataa(\my_reg[23][18]~q ),
	.datab(\Mux13~7_combout ),
	.datac(\my_reg[31][18]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux13~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~8 .lut_mask = 16'hE2CC;
defparam \Mux13~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N16
cycloneive_lcell_comb \my_reg[30][18]~feeder (
// Equation(s):
// \my_reg[30][18]~feeder_combout  = \wdat~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat15),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[30][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[30][18]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[30][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N17
dffeas \my_reg[30][18] (
	.clk(CLK),
	.d(\my_reg[30][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][18] .is_wysiwyg = "true";
defparam \my_reg[30][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N15
dffeas \my_reg[18][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][18] .is_wysiwyg = "true";
defparam \my_reg[18][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N14
cycloneive_lcell_comb \Mux13~2 (
// Equation(s):
// \Mux13~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[22][18]~q )) # (!dcifimemload_23 & ((\my_reg[18][18]~q )))))

	.dataa(\my_reg[22][18]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[18][18]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~2 .lut_mask = 16'hEE30;
defparam \Mux13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N12
cycloneive_lcell_comb \Mux13~3 (
// Equation(s):
// \Mux13~3_combout  = (dcifimemload_24 & ((\Mux13~2_combout  & ((\my_reg[30][18]~q ))) # (!\Mux13~2_combout  & (\my_reg[26][18]~q )))) # (!dcifimemload_24 & (((\Mux13~2_combout ))))

	.dataa(\my_reg[26][18]~q ),
	.datab(\my_reg[30][18]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux13~2_combout ),
	.cin(gnd),
	.combout(\Mux13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~3 .lut_mask = 16'hCFA0;
defparam \Mux13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y30_N5
dffeas \my_reg[16][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][18] .is_wysiwyg = "true";
defparam \my_reg[16][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N4
cycloneive_lcell_comb \Mux13~4 (
// Equation(s):
// \Mux13~4_combout  = (dcifimemload_23 & ((\my_reg[20][18]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[16][18]~q  & !dcifimemload_24))))

	.dataa(\my_reg[20][18]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[16][18]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~4 .lut_mask = 16'hCCB8;
defparam \Mux13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y30_N27
dffeas \my_reg[28][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][18] .is_wysiwyg = "true";
defparam \my_reg[28][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N26
cycloneive_lcell_comb \Mux13~5 (
// Equation(s):
// \Mux13~5_combout  = (\Mux13~4_combout  & (((\my_reg[28][18]~q ) # (!dcifimemload_24)))) # (!\Mux13~4_combout  & (\my_reg[24][18]~q  & ((dcifimemload_24))))

	.dataa(\my_reg[24][18]~q ),
	.datab(\Mux13~4_combout ),
	.datac(\my_reg[28][18]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux13~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~5 .lut_mask = 16'hE2CC;
defparam \Mux13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N4
cycloneive_lcell_comb \Mux13~6 (
// Equation(s):
// \Mux13~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux13~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\Mux13~5_combout ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux13~3_combout ),
	.datad(\Mux13~5_combout ),
	.cin(gnd),
	.combout(\Mux13~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~6 .lut_mask = 16'hB9A8;
defparam \Mux13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N8
cycloneive_lcell_comb \my_reg[21][18]~feeder (
// Equation(s):
// \my_reg[21][18]~feeder_combout  = \wdat~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat15),
	.cin(gnd),
	.combout(\my_reg[21][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][18]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[21][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N9
dffeas \my_reg[21][18] (
	.clk(CLK),
	.d(\my_reg[21][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][18] .is_wysiwyg = "true";
defparam \my_reg[21][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N27
dffeas \my_reg[29][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][18] .is_wysiwyg = "true";
defparam \my_reg[29][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N16
cycloneive_lcell_comb \my_reg[25][18]~feeder (
// Equation(s):
// \my_reg[25][18]~feeder_combout  = \wdat~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat15),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[25][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][18]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[25][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N17
dffeas \my_reg[25][18] (
	.clk(CLK),
	.d(\my_reg[25][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][18] .is_wysiwyg = "true";
defparam \my_reg[25][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N18
cycloneive_lcell_comb \my_reg[17][18]~feeder (
// Equation(s):
// \my_reg[17][18]~feeder_combout  = \wdat~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat15),
	.cin(gnd),
	.combout(\my_reg[17][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[17][18]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[17][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N19
dffeas \my_reg[17][18] (
	.clk(CLK),
	.d(\my_reg[17][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][18] .is_wysiwyg = "true";
defparam \my_reg[17][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N16
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (dcifimemload_24 & ((\my_reg[25][18]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((!dcifimemload_23 & \my_reg[17][18]~q ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[25][18]~q ),
	.datac(dcifimemload_23),
	.datad(\my_reg[17][18]~q ),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hADA8;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N26
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// \Mux13~1_combout  = (dcifimemload_23 & ((\Mux13~0_combout  & ((\my_reg[29][18]~q ))) # (!\Mux13~0_combout  & (\my_reg[21][18]~q )))) # (!dcifimemload_23 & (((\Mux13~0_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[21][18]~q ),
	.datac(\my_reg[29][18]~q ),
	.datad(\Mux13~0_combout ),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hF588;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N18
cycloneive_lcell_comb \Mux13~9 (
// Equation(s):
// \Mux13~9_combout  = (dcifimemload_21 & ((\Mux13~6_combout  & (\Mux13~8_combout )) # (!\Mux13~6_combout  & ((\Mux13~1_combout ))))) # (!dcifimemload_21 & (((\Mux13~6_combout ))))

	.dataa(\Mux13~8_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux13~6_combout ),
	.datad(\Mux13~1_combout ),
	.cin(gnd),
	.combout(\Mux13~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~9 .lut_mask = 16'hBCB0;
defparam \Mux13~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N22
cycloneive_lcell_comb \my_reg[13][18]~feeder (
// Equation(s):
// \my_reg[13][18]~feeder_combout  = \wdat~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat15),
	.cin(gnd),
	.combout(\my_reg[13][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[13][18]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[13][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N23
dffeas \my_reg[13][18] (
	.clk(CLK),
	.d(\my_reg[13][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][18] .is_wysiwyg = "true";
defparam \my_reg[13][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N28
cycloneive_lcell_comb \Mux45~7 (
// Equation(s):
// \Mux45~7_combout  = (dcifimemload_16 & ((\my_reg[13][18]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\my_reg[12][18]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[13][18]~q ),
	.datac(\my_reg[12][18]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux45~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~7 .lut_mask = 16'hAAD8;
defparam \Mux45~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N22
cycloneive_lcell_comb \Mux45~8 (
// Equation(s):
// \Mux45~8_combout  = (dcifimemload_17 & ((\Mux45~7_combout  & (\my_reg[15][18]~q )) # (!\Mux45~7_combout  & ((\my_reg[14][18]~q ))))) # (!dcifimemload_17 & (((\Mux45~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[15][18]~q ),
	.datac(\my_reg[14][18]~q ),
	.datad(\Mux45~7_combout ),
	.cin(gnd),
	.combout(\Mux45~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~8 .lut_mask = 16'hDDA0;
defparam \Mux45~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y30_N21
dffeas \my_reg[10][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][18] .is_wysiwyg = "true";
defparam \my_reg[10][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N20
cycloneive_lcell_comb \Mux45~0 (
// Equation(s):
// \Mux45~0_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[10][18]~q ))) # (!dcifimemload_17 & (\my_reg[8][18]~q ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[8][18]~q ),
	.datac(\my_reg[10][18]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux45~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~0 .lut_mask = 16'hFA44;
defparam \Mux45~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N22
cycloneive_lcell_comb \Mux45~1 (
// Equation(s):
// \Mux45~1_combout  = (dcifimemload_16 & ((\Mux45~0_combout  & (\my_reg[11][18]~q )) # (!\Mux45~0_combout  & ((\my_reg[9][18]~q ))))) # (!dcifimemload_16 & (((\Mux45~0_combout ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[11][18]~q ),
	.datac(\my_reg[9][18]~q ),
	.datad(\Mux45~0_combout ),
	.cin(gnd),
	.combout(\Mux45~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~1 .lut_mask = 16'hDDA0;
defparam \Mux45~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N13
dffeas \my_reg[3][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][18] .is_wysiwyg = "true";
defparam \my_reg[3][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N12
cycloneive_lcell_comb \Mux45~4 (
// Equation(s):
// \Mux45~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][18]~q ))) # (!dcifimemload_17 & (\my_reg[1][18]~q ))))

	.dataa(\my_reg[1][18]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[3][18]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux45~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~4 .lut_mask = 16'hC088;
defparam \Mux45~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N26
cycloneive_lcell_comb \Mux45~5 (
// Equation(s):
// \Mux45~5_combout  = (\Mux45~4_combout ) # ((\my_reg[2][18]~q  & (!dcifimemload_16 & dcifimemload_17)))

	.dataa(\my_reg[2][18]~q ),
	.datab(dcifimemload_16),
	.datac(dcifimemload_17),
	.datad(\Mux45~4_combout ),
	.cin(gnd),
	.combout(\Mux45~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~5 .lut_mask = 16'hFF20;
defparam \Mux45~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y32_N17
dffeas \my_reg[6][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][18] .is_wysiwyg = "true";
defparam \my_reg[6][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N16
cycloneive_lcell_comb \Mux45~3 (
// Equation(s):
// \Mux45~3_combout  = (\Mux45~2_combout  & ((\my_reg[7][18]~q ) # ((!dcifimemload_17)))) # (!\Mux45~2_combout  & (((\my_reg[6][18]~q  & dcifimemload_17))))

	.dataa(\Mux45~2_combout ),
	.datab(\my_reg[7][18]~q ),
	.datac(\my_reg[6][18]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux45~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~3 .lut_mask = 16'hD8AA;
defparam \Mux45~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N24
cycloneive_lcell_comb \Mux45~6 (
// Equation(s):
// \Mux45~6_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & ((\Mux45~3_combout ))) # (!dcifimemload_18 & (\Mux45~5_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux45~5_combout ),
	.datad(\Mux45~3_combout ),
	.cin(gnd),
	.combout(\Mux45~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~6 .lut_mask = 16'hDC98;
defparam \Mux45~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N17
dffeas \my_reg[23][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][18] .is_wysiwyg = "true";
defparam \my_reg[23][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N16
cycloneive_lcell_comb \Mux45~17 (
// Equation(s):
// \Mux45~17_combout  = (dcifimemload_18 & (((\my_reg[23][18]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[19][18]~q  & ((!dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[19][18]~q ),
	.datac(\my_reg[23][18]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux45~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~17 .lut_mask = 16'hAAE4;
defparam \Mux45~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N26
cycloneive_lcell_comb \Mux45~18 (
// Equation(s):
// \Mux45~18_combout  = (dcifimemload_19 & ((\Mux45~17_combout  & (\my_reg[31][18]~q )) # (!\Mux45~17_combout  & ((\my_reg[27][18]~q ))))) # (!dcifimemload_19 & (((\Mux45~17_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[31][18]~q ),
	.datac(\my_reg[27][18]~q ),
	.datad(\Mux45~17_combout ),
	.cin(gnd),
	.combout(\Mux45~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~18 .lut_mask = 16'hDDA0;
defparam \Mux45~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y31_N15
dffeas \my_reg[20][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][18] .is_wysiwyg = "true";
defparam \my_reg[20][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N1
dffeas \my_reg[24][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][18] .is_wysiwyg = "true";
defparam \my_reg[24][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N0
cycloneive_lcell_comb \Mux45~14 (
// Equation(s):
// \Mux45~14_combout  = (dcifimemload_19 & (((\my_reg[24][18]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[16][18]~q  & ((!dcifimemload_18))))

	.dataa(\my_reg[16][18]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[24][18]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux45~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~14 .lut_mask = 16'hCCE2;
defparam \Mux45~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N14
cycloneive_lcell_comb \Mux45~15 (
// Equation(s):
// \Mux45~15_combout  = (dcifimemload_18 & ((\Mux45~14_combout  & (\my_reg[28][18]~q )) # (!\Mux45~14_combout  & ((\my_reg[20][18]~q ))))) # (!dcifimemload_18 & (((\Mux45~14_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[28][18]~q ),
	.datac(\my_reg[20][18]~q ),
	.datad(\Mux45~14_combout ),
	.cin(gnd),
	.combout(\Mux45~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~15 .lut_mask = 16'hDDA0;
defparam \Mux45~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N6
cycloneive_lcell_comb \my_reg[22][18]~feeder (
// Equation(s):
// \my_reg[22][18]~feeder_combout  = \wdat~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat15),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[22][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[22][18]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[22][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N7
dffeas \my_reg[22][18] (
	.clk(CLK),
	.d(\my_reg[22][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][18] .is_wysiwyg = "true";
defparam \my_reg[22][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N21
dffeas \my_reg[26][18] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][18] .is_wysiwyg = "true";
defparam \my_reg[26][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N20
cycloneive_lcell_comb \Mux45~12 (
// Equation(s):
// \Mux45~12_combout  = (dcifimemload_19 & (((\my_reg[26][18]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[18][18]~q  & ((!dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[18][18]~q ),
	.datac(\my_reg[26][18]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux45~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~12 .lut_mask = 16'hAAE4;
defparam \Mux45~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N0
cycloneive_lcell_comb \Mux45~13 (
// Equation(s):
// \Mux45~13_combout  = (dcifimemload_18 & ((\Mux45~12_combout  & ((\my_reg[30][18]~q ))) # (!\Mux45~12_combout  & (\my_reg[22][18]~q )))) # (!dcifimemload_18 & (((\Mux45~12_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[22][18]~q ),
	.datac(\my_reg[30][18]~q ),
	.datad(\Mux45~12_combout ),
	.cin(gnd),
	.combout(\Mux45~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~13 .lut_mask = 16'hF588;
defparam \Mux45~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N8
cycloneive_lcell_comb \Mux45~16 (
// Equation(s):
// \Mux45~16_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux45~13_combout ))) # (!dcifimemload_17 & (\Mux45~15_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux45~15_combout ),
	.datad(\Mux45~13_combout ),
	.cin(gnd),
	.combout(\Mux45~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~16 .lut_mask = 16'hDC98;
defparam \Mux45~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N6
cycloneive_lcell_comb \Mux45~10 (
// Equation(s):
// \Mux45~10_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[21][18]~q ))) # (!dcifimemload_18 & (\my_reg[17][18]~q ))))

	.dataa(\my_reg[17][18]~q ),
	.datab(\my_reg[21][18]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux45~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~10 .lut_mask = 16'hFC0A;
defparam \Mux45~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N12
cycloneive_lcell_comb \Mux45~11 (
// Equation(s):
// \Mux45~11_combout  = (dcifimemload_19 & ((\Mux45~10_combout  & (\my_reg[29][18]~q )) # (!\Mux45~10_combout  & ((\my_reg[25][18]~q ))))) # (!dcifimemload_19 & (((\Mux45~10_combout ))))

	.dataa(\my_reg[29][18]~q ),
	.datab(\my_reg[25][18]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux45~10_combout ),
	.cin(gnd),
	.combout(\Mux45~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~11 .lut_mask = 16'hAFC0;
defparam \Mux45~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y32_N29
dffeas \my_reg[6][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][17] .is_wysiwyg = "true";
defparam \my_reg[6][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N19
dffeas \my_reg[7][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][17] .is_wysiwyg = "true";
defparam \my_reg[7][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y32_N15
dffeas \my_reg[5][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][17] .is_wysiwyg = "true";
defparam \my_reg[5][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N16
cycloneive_lcell_comb \Mux14~12 (
// Equation(s):
// \Mux14~12_combout  = (dcifimemload_21 & (((\my_reg[5][17]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\my_reg[4][17]~q  & ((!dcifimemload_22))))

	.dataa(\my_reg[4][17]~q ),
	.datab(\my_reg[5][17]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux14~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~12 .lut_mask = 16'hF0CA;
defparam \Mux14~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N18
cycloneive_lcell_comb \Mux14~13 (
// Equation(s):
// \Mux14~13_combout  = (dcifimemload_22 & ((\Mux14~12_combout  & ((\my_reg[7][17]~q ))) # (!\Mux14~12_combout  & (\my_reg[6][17]~q )))) # (!dcifimemload_22 & (((\Mux14~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[6][17]~q ),
	.datac(\my_reg[7][17]~q ),
	.datad(\Mux14~12_combout ),
	.cin(gnd),
	.combout(\Mux14~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~13 .lut_mask = 16'hF588;
defparam \Mux14~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N19
dffeas \my_reg[2][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][17] .is_wysiwyg = "true";
defparam \my_reg[2][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N23
dffeas \my_reg[1][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][17] .is_wysiwyg = "true";
defparam \my_reg[1][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N22
cycloneive_lcell_comb \Mux14~14 (
// Equation(s):
// \Mux14~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\my_reg[3][17]~q )) # (!dcifimemload_22 & ((\my_reg[1][17]~q )))))

	.dataa(\my_reg[3][17]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[1][17]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux14~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~14 .lut_mask = 16'h88C0;
defparam \Mux14~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N18
cycloneive_lcell_comb \Mux14~15 (
// Equation(s):
// \Mux14~15_combout  = (\Mux14~14_combout ) # ((!dcifimemload_21 & (dcifimemload_22 & \my_reg[2][17]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\my_reg[2][17]~q ),
	.datad(\Mux14~14_combout ),
	.cin(gnd),
	.combout(\Mux14~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~15 .lut_mask = 16'hFF40;
defparam \Mux14~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N8
cycloneive_lcell_comb \Mux14~16 (
// Equation(s):
// \Mux14~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & (\Mux14~13_combout )) # (!dcifimemload_23 & ((\Mux14~15_combout )))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux14~13_combout ),
	.datad(\Mux14~15_combout ),
	.cin(gnd),
	.combout(\Mux14~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~16 .lut_mask = 16'hD9C8;
defparam \Mux14~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N28
cycloneive_lcell_comb \my_reg[15][17]~feeder (
// Equation(s):
// \my_reg[15][17]~feeder_combout  = \wdat~33_combout 

	.dataa(wdat16),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[15][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[15][17]~feeder .lut_mask = 16'hAAAA;
defparam \my_reg[15][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N29
dffeas \my_reg[15][17] (
	.clk(CLK),
	.d(\my_reg[15][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][17] .is_wysiwyg = "true";
defparam \my_reg[15][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N7
dffeas \my_reg[14][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][17] .is_wysiwyg = "true";
defparam \my_reg[14][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N13
dffeas \my_reg[12][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][17] .is_wysiwyg = "true";
defparam \my_reg[12][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N12
cycloneive_lcell_comb \Mux14~17 (
// Equation(s):
// \Mux14~17_combout  = (dcifimemload_21 & ((\my_reg[13][17]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][17]~q  & !dcifimemload_22))))

	.dataa(\my_reg[13][17]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[12][17]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux14~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~17 .lut_mask = 16'hCCB8;
defparam \Mux14~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N6
cycloneive_lcell_comb \Mux14~18 (
// Equation(s):
// \Mux14~18_combout  = (dcifimemload_22 & ((\Mux14~17_combout  & (\my_reg[15][17]~q )) # (!\Mux14~17_combout  & ((\my_reg[14][17]~q ))))) # (!dcifimemload_22 & (((\Mux14~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[15][17]~q ),
	.datac(\my_reg[14][17]~q ),
	.datad(\Mux14~17_combout ),
	.cin(gnd),
	.combout(\Mux14~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~18 .lut_mask = 16'hDDA0;
defparam \Mux14~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N20
cycloneive_lcell_comb \my_reg[9][17]~feeder (
// Equation(s):
// \my_reg[9][17]~feeder_combout  = \wdat~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat16),
	.cin(gnd),
	.combout(\my_reg[9][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[9][17]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[9][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N21
dffeas \my_reg[9][17] (
	.clk(CLK),
	.d(\my_reg[9][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][17] .is_wysiwyg = "true";
defparam \my_reg[9][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N25
dffeas \my_reg[10][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][17] .is_wysiwyg = "true";
defparam \my_reg[10][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N24
cycloneive_lcell_comb \Mux14~10 (
// Equation(s):
// \Mux14~10_combout  = (dcifimemload_22 & (((\my_reg[10][17]~q ) # (dcifimemload_21)))) # (!dcifimemload_22 & (\my_reg[8][17]~q  & ((!dcifimemload_21))))

	.dataa(\my_reg[8][17]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[10][17]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux14~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~10 .lut_mask = 16'hCCE2;
defparam \Mux14~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N18
cycloneive_lcell_comb \Mux14~11 (
// Equation(s):
// \Mux14~11_combout  = (\Mux14~10_combout  & ((\my_reg[11][17]~q ) # ((!dcifimemload_21)))) # (!\Mux14~10_combout  & (((\my_reg[9][17]~q  & dcifimemload_21))))

	.dataa(\my_reg[11][17]~q ),
	.datab(\my_reg[9][17]~q ),
	.datac(\Mux14~10_combout ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux14~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~11 .lut_mask = 16'hACF0;
defparam \Mux14~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N14
cycloneive_lcell_comb \Mux14~19 (
// Equation(s):
// \Mux14~19_combout  = (dcifimemload_24 & ((\Mux14~16_combout  & (\Mux14~18_combout )) # (!\Mux14~16_combout  & ((\Mux14~11_combout ))))) # (!dcifimemload_24 & (\Mux14~16_combout ))

	.dataa(dcifimemload_24),
	.datab(\Mux14~16_combout ),
	.datac(\Mux14~18_combout ),
	.datad(\Mux14~11_combout ),
	.cin(gnd),
	.combout(\Mux14~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~19 .lut_mask = 16'hE6C4;
defparam \Mux14~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N29
dffeas \my_reg[27][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][17] .is_wysiwyg = "true";
defparam \my_reg[27][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y41_N3
dffeas \my_reg[31][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][17] .is_wysiwyg = "true";
defparam \my_reg[31][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y40_N31
dffeas \my_reg[23][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][17] .is_wysiwyg = "true";
defparam \my_reg[23][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y41_N1
dffeas \my_reg[19][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][17] .is_wysiwyg = "true";
defparam \my_reg[19][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N0
cycloneive_lcell_comb \Mux14~7 (
// Equation(s):
// \Mux14~7_combout  = (dcifimemload_23 & ((\my_reg[23][17]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[19][17]~q  & !dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[23][17]~q ),
	.datac(\my_reg[19][17]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux14~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~7 .lut_mask = 16'hAAD8;
defparam \Mux14~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N2
cycloneive_lcell_comb \Mux14~8 (
// Equation(s):
// \Mux14~8_combout  = (dcifimemload_24 & ((\Mux14~7_combout  & ((\my_reg[31][17]~q ))) # (!\Mux14~7_combout  & (\my_reg[27][17]~q )))) # (!dcifimemload_24 & (((\Mux14~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[27][17]~q ),
	.datac(\my_reg[31][17]~q ),
	.datad(\Mux14~7_combout ),
	.cin(gnd),
	.combout(\Mux14~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~8 .lut_mask = 16'hF588;
defparam \Mux14~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N16
cycloneive_lcell_comb \my_reg[25][17]~feeder (
// Equation(s):
// \my_reg[25][17]~feeder_combout  = \wdat~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat16),
	.cin(gnd),
	.combout(\my_reg[25][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][17]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[25][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y35_N17
dffeas \my_reg[25][17] (
	.clk(CLK),
	.d(\my_reg[25][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][17] .is_wysiwyg = "true";
defparam \my_reg[25][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N7
dffeas \my_reg[29][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][17] .is_wysiwyg = "true";
defparam \my_reg[29][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N11
dffeas \my_reg[17][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][17] .is_wysiwyg = "true";
defparam \my_reg[17][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N30
cycloneive_lcell_comb \my_reg[21][17]~feeder (
// Equation(s):
// \my_reg[21][17]~feeder_combout  = \wdat~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat16),
	.cin(gnd),
	.combout(\my_reg[21][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][17]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[21][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y35_N31
dffeas \my_reg[21][17] (
	.clk(CLK),
	.d(\my_reg[21][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][17] .is_wysiwyg = "true";
defparam \my_reg[21][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N10
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & ((\my_reg[21][17]~q ))) # (!dcifimemload_23 & (\my_reg[17][17]~q ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\my_reg[17][17]~q ),
	.datad(\my_reg[21][17]~q ),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hDC98;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N6
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// \Mux14~1_combout  = (dcifimemload_24 & ((\Mux14~0_combout  & ((\my_reg[29][17]~q ))) # (!\Mux14~0_combout  & (\my_reg[25][17]~q )))) # (!dcifimemload_24 & (((\Mux14~0_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[25][17]~q ),
	.datac(\my_reg[29][17]~q ),
	.datad(\Mux14~0_combout ),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hF588;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y30_N23
dffeas \my_reg[28][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][17] .is_wysiwyg = "true";
defparam \my_reg[28][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N29
dffeas \my_reg[16][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][17] .is_wysiwyg = "true";
defparam \my_reg[16][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N28
cycloneive_lcell_comb \Mux14~4 (
// Equation(s):
// \Mux14~4_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[24][17]~q )) # (!dcifimemload_24 & ((\my_reg[16][17]~q )))))

	.dataa(\my_reg[24][17]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[16][17]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux14~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~4 .lut_mask = 16'hEE30;
defparam \Mux14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N22
cycloneive_lcell_comb \Mux14~5 (
// Equation(s):
// \Mux14~5_combout  = (dcifimemload_23 & ((\Mux14~4_combout  & ((\my_reg[28][17]~q ))) # (!\Mux14~4_combout  & (\my_reg[20][17]~q )))) # (!dcifimemload_23 & (((\Mux14~4_combout ))))

	.dataa(\my_reg[20][17]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[28][17]~q ),
	.datad(\Mux14~4_combout ),
	.cin(gnd),
	.combout(\Mux14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~5 .lut_mask = 16'hF388;
defparam \Mux14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y42_N29
dffeas \my_reg[22][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][17] .is_wysiwyg = "true";
defparam \my_reg[22][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y42_N29
dffeas \my_reg[30][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][17] .is_wysiwyg = "true";
defparam \my_reg[30][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N0
cycloneive_lcell_comb \my_reg[18][17]~feeder (
// Equation(s):
// \my_reg[18][17]~feeder_combout  = \wdat~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat16),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[18][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[18][17]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[18][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N1
dffeas \my_reg[18][17] (
	.clk(CLK),
	.d(\my_reg[18][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][17] .is_wysiwyg = "true";
defparam \my_reg[18][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N18
cycloneive_lcell_comb \Mux14~2 (
// Equation(s):
// \Mux14~2_combout  = (dcifimemload_24 & ((\my_reg[26][17]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\my_reg[18][17]~q  & !dcifimemload_23))))

	.dataa(\my_reg[26][17]~q ),
	.datab(\my_reg[18][17]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux14~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~2 .lut_mask = 16'hF0AC;
defparam \Mux14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N28
cycloneive_lcell_comb \Mux14~3 (
// Equation(s):
// \Mux14~3_combout  = (dcifimemload_23 & ((\Mux14~2_combout  & ((\my_reg[30][17]~q ))) # (!\Mux14~2_combout  & (\my_reg[22][17]~q )))) # (!dcifimemload_23 & (((\Mux14~2_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[22][17]~q ),
	.datac(\my_reg[30][17]~q ),
	.datad(\Mux14~2_combout ),
	.cin(gnd),
	.combout(\Mux14~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~3 .lut_mask = 16'hF588;
defparam \Mux14~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N14
cycloneive_lcell_comb \Mux14~6 (
// Equation(s):
// \Mux14~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux14~3_combout ))) # (!dcifimemload_22 & (\Mux14~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux14~5_combout ),
	.datad(\Mux14~3_combout ),
	.cin(gnd),
	.combout(\Mux14~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~6 .lut_mask = 16'hDC98;
defparam \Mux14~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N10
cycloneive_lcell_comb \Mux14~9 (
// Equation(s):
// \Mux14~9_combout  = (dcifimemload_21 & ((\Mux14~6_combout  & (\Mux14~8_combout )) # (!\Mux14~6_combout  & ((\Mux14~1_combout ))))) # (!dcifimemload_21 & (((\Mux14~6_combout ))))

	.dataa(\Mux14~8_combout ),
	.datab(\Mux14~1_combout ),
	.datac(dcifimemload_21),
	.datad(\Mux14~6_combout ),
	.cin(gnd),
	.combout(\Mux14~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~9 .lut_mask = 16'hAFC0;
defparam \Mux14~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N26
cycloneive_lcell_comb \my_reg[4][17]~feeder (
// Equation(s):
// \my_reg[4][17]~feeder_combout  = \wdat~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat16),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[4][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[4][17]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[4][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y42_N27
dffeas \my_reg[4][17] (
	.clk(CLK),
	.d(\my_reg[4][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][17] .is_wysiwyg = "true";
defparam \my_reg[4][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N14
cycloneive_lcell_comb \Mux46~0 (
// Equation(s):
// \Mux46~0_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][17]~q ))) # (!dcifimemload_16 & (\my_reg[4][17]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[4][17]~q ),
	.datac(\my_reg[5][17]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux46~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~0 .lut_mask = 16'hFA44;
defparam \Mux46~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N28
cycloneive_lcell_comb \Mux46~1 (
// Equation(s):
// \Mux46~1_combout  = (\Mux46~0_combout  & ((\my_reg[7][17]~q ) # ((!dcifimemload_17)))) # (!\Mux46~0_combout  & (((\my_reg[6][17]~q  & dcifimemload_17))))

	.dataa(\my_reg[7][17]~q ),
	.datab(\Mux46~0_combout ),
	.datac(\my_reg[6][17]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux46~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~1 .lut_mask = 16'hB8CC;
defparam \Mux46~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N26
cycloneive_lcell_comb \my_reg[13][17]~feeder (
// Equation(s):
// \my_reg[13][17]~feeder_combout  = \wdat~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat16),
	.cin(gnd),
	.combout(\my_reg[13][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[13][17]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[13][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y31_N27
dffeas \my_reg[13][17] (
	.clk(CLK),
	.d(\my_reg[13][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][17] .is_wysiwyg = "true";
defparam \my_reg[13][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N4
cycloneive_lcell_comb \Mux46~7 (
// Equation(s):
// \Mux46~7_combout  = (dcifimemload_16 & (((\my_reg[13][17]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[12][17]~q  & ((!dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[12][17]~q ),
	.datac(\my_reg[13][17]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux46~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~7 .lut_mask = 16'hAAE4;
defparam \Mux46~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N26
cycloneive_lcell_comb \Mux46~8 (
// Equation(s):
// \Mux46~8_combout  = (dcifimemload_17 & ((\Mux46~7_combout  & (\my_reg[15][17]~q )) # (!\Mux46~7_combout  & ((\my_reg[14][17]~q ))))) # (!dcifimemload_17 & (((\Mux46~7_combout ))))

	.dataa(\my_reg[15][17]~q ),
	.datab(\my_reg[14][17]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux46~7_combout ),
	.cin(gnd),
	.combout(\Mux46~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~8 .lut_mask = 16'hAFC0;
defparam \Mux46~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N25
dffeas \my_reg[3][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][17] .is_wysiwyg = "true";
defparam \my_reg[3][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N24
cycloneive_lcell_comb \Mux46~4 (
// Equation(s):
// \Mux46~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][17]~q ))) # (!dcifimemload_17 & (\my_reg[1][17]~q ))))

	.dataa(\my_reg[1][17]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[3][17]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux46~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~4 .lut_mask = 16'hC088;
defparam \Mux46~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N22
cycloneive_lcell_comb \Mux46~5 (
// Equation(s):
// \Mux46~5_combout  = (\Mux46~4_combout ) # ((\my_reg[2][17]~q  & (!dcifimemload_16 & dcifimemload_17)))

	.dataa(\my_reg[2][17]~q ),
	.datab(dcifimemload_16),
	.datac(dcifimemload_17),
	.datad(\Mux46~4_combout ),
	.cin(gnd),
	.combout(\Mux46~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~5 .lut_mask = 16'hFF20;
defparam \Mux46~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N5
dffeas \my_reg[8][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][17] .is_wysiwyg = "true";
defparam \my_reg[8][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N4
cycloneive_lcell_comb \Mux46~2 (
// Equation(s):
// \Mux46~2_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\my_reg[10][17]~q )) # (!dcifimemload_17 & ((\my_reg[8][17]~q )))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[10][17]~q ),
	.datac(\my_reg[8][17]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux46~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~2 .lut_mask = 16'hEE50;
defparam \Mux46~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N7
dffeas \my_reg[11][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][17] .is_wysiwyg = "true";
defparam \my_reg[11][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N6
cycloneive_lcell_comb \Mux46~3 (
// Equation(s):
// \Mux46~3_combout  = (\Mux46~2_combout  & (((\my_reg[11][17]~q ) # (!dcifimemload_16)))) # (!\Mux46~2_combout  & (\my_reg[9][17]~q  & ((dcifimemload_16))))

	.dataa(\my_reg[9][17]~q ),
	.datab(\Mux46~2_combout ),
	.datac(\my_reg[11][17]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux46~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~3 .lut_mask = 16'hE2CC;
defparam \Mux46~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N28
cycloneive_lcell_comb \Mux46~6 (
// Equation(s):
// \Mux46~6_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & ((\Mux46~3_combout ))) # (!dcifimemload_19 & (\Mux46~5_combout ))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux46~5_combout ),
	.datad(\Mux46~3_combout ),
	.cin(gnd),
	.combout(\Mux46~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~6 .lut_mask = 16'hDC98;
defparam \Mux46~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N24
cycloneive_lcell_comb \Mux46~10 (
// Equation(s):
// \Mux46~10_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[25][17]~q ))) # (!dcifimemload_19 & (\my_reg[17][17]~q ))))

	.dataa(\my_reg[17][17]~q ),
	.datab(\my_reg[25][17]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux46~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~10 .lut_mask = 16'hFC0A;
defparam \Mux46~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N10
cycloneive_lcell_comb \Mux46~11 (
// Equation(s):
// \Mux46~11_combout  = (dcifimemload_18 & ((\Mux46~10_combout  & ((\my_reg[29][17]~q ))) # (!\Mux46~10_combout  & (\my_reg[21][17]~q )))) # (!dcifimemload_18 & (((\Mux46~10_combout ))))

	.dataa(\my_reg[21][17]~q ),
	.datab(\my_reg[29][17]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux46~10_combout ),
	.cin(gnd),
	.combout(\Mux46~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~11 .lut_mask = 16'hCFA0;
defparam \Mux46~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N28
cycloneive_lcell_comb \Mux46~17 (
// Equation(s):
// \Mux46~17_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[27][17]~q ))) # (!dcifimemload_19 & (\my_reg[19][17]~q ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[19][17]~q ),
	.datac(\my_reg[27][17]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux46~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~17 .lut_mask = 16'hFA44;
defparam \Mux46~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N30
cycloneive_lcell_comb \Mux46~18 (
// Equation(s):
// \Mux46~18_combout  = (dcifimemload_18 & ((\Mux46~17_combout  & (\my_reg[31][17]~q )) # (!\Mux46~17_combout  & ((\my_reg[23][17]~q ))))) # (!dcifimemload_18 & (((\Mux46~17_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[31][17]~q ),
	.datac(\my_reg[23][17]~q ),
	.datad(\Mux46~17_combout ),
	.cin(gnd),
	.combout(\Mux46~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~18 .lut_mask = 16'hDDA0;
defparam \Mux46~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N8
cycloneive_lcell_comb \my_reg[24][17]~feeder (
// Equation(s):
// \my_reg[24][17]~feeder_combout  = \wdat~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat16),
	.cin(gnd),
	.combout(\my_reg[24][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[24][17]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[24][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y31_N9
dffeas \my_reg[24][17] (
	.clk(CLK),
	.d(\my_reg[24][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][17] .is_wysiwyg = "true";
defparam \my_reg[24][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N6
cycloneive_lcell_comb \Mux46~14 (
// Equation(s):
// \Mux46~14_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\my_reg[20][17]~q )) # (!dcifimemload_18 & ((\my_reg[16][17]~q )))))

	.dataa(\my_reg[20][17]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[16][17]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux46~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~14 .lut_mask = 16'hEE30;
defparam \Mux46~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N4
cycloneive_lcell_comb \Mux46~15 (
// Equation(s):
// \Mux46~15_combout  = (dcifimemload_19 & ((\Mux46~14_combout  & (\my_reg[28][17]~q )) # (!\Mux46~14_combout  & ((\my_reg[24][17]~q ))))) # (!dcifimemload_19 & (((\Mux46~14_combout ))))

	.dataa(\my_reg[28][17]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[24][17]~q ),
	.datad(\Mux46~14_combout ),
	.cin(gnd),
	.combout(\Mux46~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~15 .lut_mask = 16'hBBC0;
defparam \Mux46~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y42_N23
dffeas \my_reg[26][17] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][17] .is_wysiwyg = "true";
defparam \my_reg[26][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N28
cycloneive_lcell_comb \Mux46~12 (
// Equation(s):
// \Mux46~12_combout  = (dcifimemload_18 & (((\my_reg[22][17]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[18][17]~q  & ((!dcifimemload_19))))

	.dataa(\my_reg[18][17]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[22][17]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux46~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~12 .lut_mask = 16'hCCE2;
defparam \Mux46~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N22
cycloneive_lcell_comb \Mux46~13 (
// Equation(s):
// \Mux46~13_combout  = (dcifimemload_19 & ((\Mux46~12_combout  & (\my_reg[30][17]~q )) # (!\Mux46~12_combout  & ((\my_reg[26][17]~q ))))) # (!dcifimemload_19 & (((\Mux46~12_combout ))))

	.dataa(\my_reg[30][17]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[26][17]~q ),
	.datad(\Mux46~12_combout ),
	.cin(gnd),
	.combout(\Mux46~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~13 .lut_mask = 16'hBBC0;
defparam \Mux46~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N10
cycloneive_lcell_comb \Mux46~16 (
// Equation(s):
// \Mux46~16_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux46~13_combout ))) # (!dcifimemload_17 & (\Mux46~15_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux46~15_combout ),
	.datad(\Mux46~13_combout ),
	.cin(gnd),
	.combout(\Mux46~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~16 .lut_mask = 16'hDC98;
defparam \Mux46~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N19
dffeas \my_reg[2][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][16] .is_wysiwyg = "true";
defparam \my_reg[2][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N25
dffeas \my_reg[1][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][16] .is_wysiwyg = "true";
defparam \my_reg[1][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y42_N19
dffeas \my_reg[3][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][16] .is_wysiwyg = "true";
defparam \my_reg[3][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N24
cycloneive_lcell_comb \Mux15~14 (
// Equation(s):
// \Mux15~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][16]~q ))) # (!dcifimemload_22 & (\my_reg[1][16]~q ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\my_reg[1][16]~q ),
	.datad(\my_reg[3][16]~q ),
	.cin(gnd),
	.combout(\Mux15~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~14 .lut_mask = 16'hA820;
defparam \Mux15~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N18
cycloneive_lcell_comb \Mux15~15 (
// Equation(s):
// \Mux15~15_combout  = (\Mux15~14_combout ) # ((!dcifimemload_21 & (dcifimemload_22 & \my_reg[2][16]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\my_reg[2][16]~q ),
	.datad(\Mux15~14_combout ),
	.cin(gnd),
	.combout(\Mux15~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~15 .lut_mask = 16'hFF40;
defparam \Mux15~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y30_N7
dffeas \my_reg[9][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][16] .is_wysiwyg = "true";
defparam \my_reg[9][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y41_N31
dffeas \my_reg[11][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][16] .is_wysiwyg = "true";
defparam \my_reg[11][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N17
dffeas \my_reg[10][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][16] .is_wysiwyg = "true";
defparam \my_reg[10][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y41_N29
dffeas \my_reg[8][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][16] .is_wysiwyg = "true";
defparam \my_reg[8][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N28
cycloneive_lcell_comb \Mux15~12 (
// Equation(s):
// \Mux15~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][16]~q )) # (!dcifimemload_22 & ((\my_reg[8][16]~q )))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[10][16]~q ),
	.datac(\my_reg[8][16]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux15~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~12 .lut_mask = 16'hEE50;
defparam \Mux15~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N30
cycloneive_lcell_comb \Mux15~13 (
// Equation(s):
// \Mux15~13_combout  = (dcifimemload_21 & ((\Mux15~12_combout  & ((\my_reg[11][16]~q ))) # (!\Mux15~12_combout  & (\my_reg[9][16]~q )))) # (!dcifimemload_21 & (((\Mux15~12_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][16]~q ),
	.datac(\my_reg[11][16]~q ),
	.datad(\Mux15~12_combout ),
	.cin(gnd),
	.combout(\Mux15~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~13 .lut_mask = 16'hF588;
defparam \Mux15~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N20
cycloneive_lcell_comb \Mux15~16 (
// Equation(s):
// \Mux15~16_combout  = (dcifimemload_24 & (((dcifimemload_23) # (\Mux15~13_combout )))) # (!dcifimemload_24 & (\Mux15~15_combout  & (!dcifimemload_23)))

	.dataa(dcifimemload_24),
	.datab(\Mux15~15_combout ),
	.datac(dcifimemload_23),
	.datad(\Mux15~13_combout ),
	.cin(gnd),
	.combout(\Mux15~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~16 .lut_mask = 16'hAEA4;
defparam \Mux15~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N21
dffeas \my_reg[14][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][16] .is_wysiwyg = "true";
defparam \my_reg[14][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N15
dffeas \my_reg[15][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][16] .is_wysiwyg = "true";
defparam \my_reg[15][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N15
dffeas \my_reg[12][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][16] .is_wysiwyg = "true";
defparam \my_reg[12][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N14
cycloneive_lcell_comb \Mux15~17 (
// Equation(s):
// \Mux15~17_combout  = (dcifimemload_21 & ((\my_reg[13][16]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][16]~q  & !dcifimemload_22))))

	.dataa(\my_reg[13][16]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[12][16]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux15~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~17 .lut_mask = 16'hCCB8;
defparam \Mux15~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N14
cycloneive_lcell_comb \Mux15~18 (
// Equation(s):
// \Mux15~18_combout  = (dcifimemload_22 & ((\Mux15~17_combout  & ((\my_reg[15][16]~q ))) # (!\Mux15~17_combout  & (\my_reg[14][16]~q )))) # (!dcifimemload_22 & (((\Mux15~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[14][16]~q ),
	.datac(\my_reg[15][16]~q ),
	.datad(\Mux15~17_combout ),
	.cin(gnd),
	.combout(\Mux15~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~18 .lut_mask = 16'hF588;
defparam \Mux15~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N23
dffeas \my_reg[7][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][16] .is_wysiwyg = "true";
defparam \my_reg[7][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N15
dffeas \my_reg[6][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][16] .is_wysiwyg = "true";
defparam \my_reg[6][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N9
dffeas \my_reg[4][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][16] .is_wysiwyg = "true";
defparam \my_reg[4][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N25
dffeas \my_reg[5][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][16] .is_wysiwyg = "true";
defparam \my_reg[5][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N24
cycloneive_lcell_comb \Mux15~10 (
// Equation(s):
// \Mux15~10_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\my_reg[5][16]~q ))) # (!dcifimemload_21 & (\my_reg[4][16]~q ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[4][16]~q ),
	.datac(\my_reg[5][16]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux15~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~10 .lut_mask = 16'hFA44;
defparam \Mux15~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N14
cycloneive_lcell_comb \Mux15~11 (
// Equation(s):
// \Mux15~11_combout  = (dcifimemload_22 & ((\Mux15~10_combout  & (\my_reg[7][16]~q )) # (!\Mux15~10_combout  & ((\my_reg[6][16]~q ))))) # (!dcifimemload_22 & (((\Mux15~10_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[7][16]~q ),
	.datac(\my_reg[6][16]~q ),
	.datad(\Mux15~10_combout ),
	.cin(gnd),
	.combout(\Mux15~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~11 .lut_mask = 16'hDDA0;
defparam \Mux15~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N14
cycloneive_lcell_comb \Mux15~19 (
// Equation(s):
// \Mux15~19_combout  = (dcifimemload_23 & ((\Mux15~16_combout  & (\Mux15~18_combout )) # (!\Mux15~16_combout  & ((\Mux15~11_combout ))))) # (!dcifimemload_23 & (\Mux15~16_combout ))

	.dataa(dcifimemload_23),
	.datab(\Mux15~16_combout ),
	.datac(\Mux15~18_combout ),
	.datad(\Mux15~11_combout ),
	.cin(gnd),
	.combout(\Mux15~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~19 .lut_mask = 16'hE6C4;
defparam \Mux15~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N26
cycloneive_lcell_comb \my_reg[23][16]~feeder (
// Equation(s):
// \my_reg[23][16]~feeder_combout  = \wdat~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat17),
	.cin(gnd),
	.combout(\my_reg[23][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[23][16]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[23][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N27
dffeas \my_reg[23][16] (
	.clk(CLK),
	.d(\my_reg[23][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][16] .is_wysiwyg = "true";
defparam \my_reg[23][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y41_N31
dffeas \my_reg[31][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][16] .is_wysiwyg = "true";
defparam \my_reg[31][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N28
cycloneive_lcell_comb \my_reg[27][16]~feeder (
// Equation(s):
// \my_reg[27][16]~feeder_combout  = \wdat~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat17),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[27][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[27][16]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[27][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N29
dffeas \my_reg[27][16] (
	.clk(CLK),
	.d(\my_reg[27][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][16] .is_wysiwyg = "true";
defparam \my_reg[27][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y41_N13
dffeas \my_reg[19][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][16] .is_wysiwyg = "true";
defparam \my_reg[19][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N12
cycloneive_lcell_comb \Mux15~7 (
// Equation(s):
// \Mux15~7_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[27][16]~q )) # (!dcifimemload_24 & ((\my_reg[19][16]~q )))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[27][16]~q ),
	.datac(\my_reg[19][16]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux15~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~7 .lut_mask = 16'hEE50;
defparam \Mux15~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N30
cycloneive_lcell_comb \Mux15~8 (
// Equation(s):
// \Mux15~8_combout  = (dcifimemload_23 & ((\Mux15~7_combout  & ((\my_reg[31][16]~q ))) # (!\Mux15~7_combout  & (\my_reg[23][16]~q )))) # (!dcifimemload_23 & (((\Mux15~7_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[23][16]~q ),
	.datac(\my_reg[31][16]~q ),
	.datad(\Mux15~7_combout ),
	.cin(gnd),
	.combout(\Mux15~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~8 .lut_mask = 16'hF588;
defparam \Mux15~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N17
dffeas \my_reg[29][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][16] .is_wysiwyg = "true";
defparam \my_reg[29][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N6
cycloneive_lcell_comb \my_reg[25][16]~feeder (
// Equation(s):
// \my_reg[25][16]~feeder_combout  = \wdat~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat17),
	.cin(gnd),
	.combout(\my_reg[25][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][16]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[25][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N7
dffeas \my_reg[25][16] (
	.clk(CLK),
	.d(\my_reg[25][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][16] .is_wysiwyg = "true";
defparam \my_reg[25][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N17
dffeas \my_reg[17][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][16] .is_wysiwyg = "true";
defparam \my_reg[17][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N16
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[25][16]~q )) # (!dcifimemload_24 & ((\my_reg[17][16]~q )))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[25][16]~q ),
	.datac(\my_reg[17][16]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hEE50;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N16
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// \Mux15~1_combout  = (dcifimemload_23 & ((\Mux15~0_combout  & ((\my_reg[29][16]~q ))) # (!\Mux15~0_combout  & (\my_reg[21][16]~q )))) # (!dcifimemload_23 & (((\Mux15~0_combout ))))

	.dataa(\my_reg[21][16]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[29][16]~q ),
	.datad(\Mux15~0_combout ),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hF388;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N30
cycloneive_lcell_comb \my_reg[24][16]~feeder (
// Equation(s):
// \my_reg[24][16]~feeder_combout  = \wdat~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat17),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[24][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[24][16]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[24][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N31
dffeas \my_reg[24][16] (
	.clk(CLK),
	.d(\my_reg[24][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][16] .is_wysiwyg = "true";
defparam \my_reg[24][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N13
dffeas \my_reg[28][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][16] .is_wysiwyg = "true";
defparam \my_reg[28][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N20
cycloneive_lcell_comb \my_reg[16][16]~feeder (
// Equation(s):
// \my_reg[16][16]~feeder_combout  = \wdat~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat17),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[16][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[16][16]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[16][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N21
dffeas \my_reg[16][16] (
	.clk(CLK),
	.d(\my_reg[16][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][16] .is_wysiwyg = "true";
defparam \my_reg[16][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N22
cycloneive_lcell_comb \Mux15~4 (
// Equation(s):
// \Mux15~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[20][16]~q )) # (!dcifimemload_23 & ((\my_reg[16][16]~q )))))

	.dataa(\my_reg[20][16]~q ),
	.datab(\my_reg[16][16]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux15~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~4 .lut_mask = 16'hFA0C;
defparam \Mux15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N12
cycloneive_lcell_comb \Mux15~5 (
// Equation(s):
// \Mux15~5_combout  = (dcifimemload_24 & ((\Mux15~4_combout  & ((\my_reg[28][16]~q ))) # (!\Mux15~4_combout  & (\my_reg[24][16]~q )))) # (!dcifimemload_24 & (((\Mux15~4_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[24][16]~q ),
	.datac(\my_reg[28][16]~q ),
	.datad(\Mux15~4_combout ),
	.cin(gnd),
	.combout(\Mux15~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~5 .lut_mask = 16'hF588;
defparam \Mux15~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N0
cycloneive_lcell_comb \Mux15~6 (
// Equation(s):
// \Mux15~6_combout  = (dcifimemload_22 & ((\Mux15~3_combout ) # ((dcifimemload_21)))) # (!dcifimemload_22 & (((!dcifimemload_21 & \Mux15~5_combout ))))

	.dataa(\Mux15~3_combout ),
	.datab(dcifimemload_22),
	.datac(dcifimemload_21),
	.datad(\Mux15~5_combout ),
	.cin(gnd),
	.combout(\Mux15~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~6 .lut_mask = 16'hCBC8;
defparam \Mux15~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N2
cycloneive_lcell_comb \Mux15~9 (
// Equation(s):
// \Mux15~9_combout  = (dcifimemload_21 & ((\Mux15~6_combout  & (\Mux15~8_combout )) # (!\Mux15~6_combout  & ((\Mux15~1_combout ))))) # (!dcifimemload_21 & (((\Mux15~6_combout ))))

	.dataa(\Mux15~8_combout ),
	.datab(\Mux15~1_combout ),
	.datac(dcifimemload_21),
	.datad(\Mux15~6_combout ),
	.cin(gnd),
	.combout(\Mux15~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~9 .lut_mask = 16'hAFC0;
defparam \Mux15~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N16
cycloneive_lcell_comb \Mux47~0 (
// Equation(s):
// \Mux47~0_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[10][16]~q ))) # (!dcifimemload_17 & (\my_reg[8][16]~q ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[8][16]~q ),
	.datac(\my_reg[10][16]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux47~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~0 .lut_mask = 16'hFA44;
defparam \Mux47~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N6
cycloneive_lcell_comb \Mux47~1 (
// Equation(s):
// \Mux47~1_combout  = (\Mux47~0_combout  & ((\my_reg[11][16]~q ) # ((!dcifimemload_16)))) # (!\Mux47~0_combout  & (((\my_reg[9][16]~q  & dcifimemload_16))))

	.dataa(\my_reg[11][16]~q ),
	.datab(\Mux47~0_combout ),
	.datac(\my_reg[9][16]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux47~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~1 .lut_mask = 16'hB8CC;
defparam \Mux47~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N9
dffeas \my_reg[13][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][16] .is_wysiwyg = "true";
defparam \my_reg[13][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N8
cycloneive_lcell_comb \Mux47~7 (
// Equation(s):
// \Mux47~7_combout  = (dcifimemload_16 & (((\my_reg[13][16]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[12][16]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[12][16]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[13][16]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux47~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~7 .lut_mask = 16'hCCE2;
defparam \Mux47~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N20
cycloneive_lcell_comb \Mux47~8 (
// Equation(s):
// \Mux47~8_combout  = (dcifimemload_17 & ((\Mux47~7_combout  & (\my_reg[15][16]~q )) # (!\Mux47~7_combout  & ((\my_reg[14][16]~q ))))) # (!dcifimemload_17 & (((\Mux47~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[15][16]~q ),
	.datac(\my_reg[14][16]~q ),
	.datad(\Mux47~7_combout ),
	.cin(gnd),
	.combout(\Mux47~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~8 .lut_mask = 16'hDDA0;
defparam \Mux47~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N8
cycloneive_lcell_comb \Mux47~2 (
// Equation(s):
// \Mux47~2_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\my_reg[5][16]~q )) # (!dcifimemload_16 & ((\my_reg[4][16]~q )))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[5][16]~q ),
	.datac(\my_reg[4][16]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux47~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~2 .lut_mask = 16'hEE50;
defparam \Mux47~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N22
cycloneive_lcell_comb \Mux47~3 (
// Equation(s):
// \Mux47~3_combout  = (\Mux47~2_combout  & (((\my_reg[7][16]~q ) # (!dcifimemload_17)))) # (!\Mux47~2_combout  & (\my_reg[6][16]~q  & ((dcifimemload_17))))

	.dataa(\my_reg[6][16]~q ),
	.datab(\Mux47~2_combout ),
	.datac(\my_reg[7][16]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux47~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~3 .lut_mask = 16'hE2CC;
defparam \Mux47~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N18
cycloneive_lcell_comb \Mux47~4 (
// Equation(s):
// \Mux47~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][16]~q ))) # (!dcifimemload_17 & (\my_reg[1][16]~q ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[1][16]~q ),
	.datac(\my_reg[3][16]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux47~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~4 .lut_mask = 16'hA088;
defparam \Mux47~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N4
cycloneive_lcell_comb \Mux47~5 (
// Equation(s):
// \Mux47~5_combout  = (\Mux47~4_combout ) # ((!dcifimemload_16 & (\my_reg[2][16]~q  & dcifimemload_17)))

	.dataa(dcifimemload_16),
	.datab(\my_reg[2][16]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux47~4_combout ),
	.cin(gnd),
	.combout(\Mux47~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~5 .lut_mask = 16'hFF40;
defparam \Mux47~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N18
cycloneive_lcell_comb \Mux47~6 (
// Equation(s):
// \Mux47~6_combout  = (dcifimemload_18 & ((dcifimemload_19) # ((\Mux47~3_combout )))) # (!dcifimemload_18 & (!dcifimemload_19 & ((\Mux47~5_combout ))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux47~3_combout ),
	.datad(\Mux47~5_combout ),
	.cin(gnd),
	.combout(\Mux47~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~6 .lut_mask = 16'hB9A8;
defparam \Mux47~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N27
dffeas \my_reg[21][16] (
	.clk(CLK),
	.d(wdat17),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][16] .is_wysiwyg = "true";
defparam \my_reg[21][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N4
cycloneive_lcell_comb \Mux47~10 (
// Equation(s):
// \Mux47~10_combout  = (dcifimemload_18 & (((\my_reg[21][16]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[17][16]~q  & ((!dcifimemload_19))))

	.dataa(\my_reg[17][16]~q ),
	.datab(\my_reg[21][16]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux47~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~10 .lut_mask = 16'hF0CA;
defparam \Mux47~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N30
cycloneive_lcell_comb \Mux47~11 (
// Equation(s):
// \Mux47~11_combout  = (\Mux47~10_combout  & (((\my_reg[29][16]~q ) # (!dcifimemload_19)))) # (!\Mux47~10_combout  & (\my_reg[25][16]~q  & ((dcifimemload_19))))

	.dataa(\my_reg[25][16]~q ),
	.datab(\Mux47~10_combout ),
	.datac(\my_reg[29][16]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux47~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~11 .lut_mask = 16'hE2CC;
defparam \Mux47~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y30_N17
dffeas \my_reg[22][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][16] .is_wysiwyg = "true";
defparam \my_reg[22][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N9
dffeas \my_reg[18][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][16] .is_wysiwyg = "true";
defparam \my_reg[18][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N27
dffeas \my_reg[26][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][16] .is_wysiwyg = "true";
defparam \my_reg[26][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N26
cycloneive_lcell_comb \Mux47~12 (
// Equation(s):
// \Mux47~12_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[26][16]~q ))) # (!dcifimemload_19 & (\my_reg[18][16]~q ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[18][16]~q ),
	.datac(\my_reg[26][16]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux47~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~12 .lut_mask = 16'hFA44;
defparam \Mux47~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N16
cycloneive_lcell_comb \Mux47~13 (
// Equation(s):
// \Mux47~13_combout  = (dcifimemload_18 & ((\Mux47~12_combout  & (\my_reg[30][16]~q )) # (!\Mux47~12_combout  & ((\my_reg[22][16]~q ))))) # (!dcifimemload_18 & (((\Mux47~12_combout ))))

	.dataa(\my_reg[30][16]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[22][16]~q ),
	.datad(\Mux47~12_combout ),
	.cin(gnd),
	.combout(\Mux47~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~13 .lut_mask = 16'hBBC0;
defparam \Mux47~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y30_N11
dffeas \my_reg[20][16] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][16] .is_wysiwyg = "true";
defparam \my_reg[20][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N8
cycloneive_lcell_comb \Mux47~14 (
// Equation(s):
// \Mux47~14_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\my_reg[24][16]~q )) # (!dcifimemload_19 & ((\my_reg[16][16]~q )))))

	.dataa(\my_reg[24][16]~q ),
	.datab(\my_reg[16][16]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux47~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~14 .lut_mask = 16'hFA0C;
defparam \Mux47~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N10
cycloneive_lcell_comb \Mux47~15 (
// Equation(s):
// \Mux47~15_combout  = (dcifimemload_18 & ((\Mux47~14_combout  & (\my_reg[28][16]~q )) # (!\Mux47~14_combout  & ((\my_reg[20][16]~q ))))) # (!dcifimemload_18 & (((\Mux47~14_combout ))))

	.dataa(\my_reg[28][16]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[20][16]~q ),
	.datad(\Mux47~14_combout ),
	.cin(gnd),
	.combout(\Mux47~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~15 .lut_mask = 16'hBBC0;
defparam \Mux47~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N8
cycloneive_lcell_comb \Mux47~16 (
// Equation(s):
// \Mux47~16_combout  = (dcifimemload_17 & ((\Mux47~13_combout ) # ((dcifimemload_16)))) # (!dcifimemload_17 & (((!dcifimemload_16 & \Mux47~15_combout ))))

	.dataa(dcifimemload_17),
	.datab(\Mux47~13_combout ),
	.datac(dcifimemload_16),
	.datad(\Mux47~15_combout ),
	.cin(gnd),
	.combout(\Mux47~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~16 .lut_mask = 16'hADA8;
defparam \Mux47~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N12
cycloneive_lcell_comb \Mux47~17 (
// Equation(s):
// \Mux47~17_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\my_reg[23][16]~q )) # (!dcifimemload_18 & ((\my_reg[19][16]~q )))))

	.dataa(\my_reg[23][16]~q ),
	.datab(\my_reg[19][16]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux47~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~17 .lut_mask = 16'hFA0C;
defparam \Mux47~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N22
cycloneive_lcell_comb \Mux47~18 (
// Equation(s):
// \Mux47~18_combout  = (dcifimemload_19 & ((\Mux47~17_combout  & (\my_reg[31][16]~q )) # (!\Mux47~17_combout  & ((\my_reg[27][16]~q ))))) # (!dcifimemload_19 & (((\Mux47~17_combout ))))

	.dataa(\my_reg[31][16]~q ),
	.datab(\my_reg[27][16]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux47~17_combout ),
	.cin(gnd),
	.combout(\Mux47~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~18 .lut_mask = 16'hAFC0;
defparam \Mux47~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N17
dffeas \my_reg[19][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][15] .is_wysiwyg = "true";
defparam \my_reg[19][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N16
cycloneive_lcell_comb \Mux16~7 (
// Equation(s):
// \Mux16~7_combout  = (dcifimemload_23 & ((\my_reg[23][15]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[19][15]~q  & !dcifimemload_24))))

	.dataa(\my_reg[23][15]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[19][15]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux16~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~7 .lut_mask = 16'hCCB8;
defparam \Mux16~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N15
dffeas \my_reg[31][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][15] .is_wysiwyg = "true";
defparam \my_reg[31][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N14
cycloneive_lcell_comb \Mux16~8 (
// Equation(s):
// \Mux16~8_combout  = (\Mux16~7_combout  & (((\my_reg[31][15]~q ) # (!dcifimemload_24)))) # (!\Mux16~7_combout  & (\my_reg[27][15]~q  & ((dcifimemload_24))))

	.dataa(\my_reg[27][15]~q ),
	.datab(\Mux16~7_combout ),
	.datac(\my_reg[31][15]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux16~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~8 .lut_mask = 16'hE2CC;
defparam \Mux16~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N21
dffeas \my_reg[22][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][15] .is_wysiwyg = "true";
defparam \my_reg[22][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N10
cycloneive_lcell_comb \my_reg[30][15]~feeder (
// Equation(s):
// \my_reg[30][15]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat18),
	.cin(gnd),
	.combout(\my_reg[30][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[30][15]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[30][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y42_N11
dffeas \my_reg[30][15] (
	.clk(CLK),
	.d(\my_reg[30][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][15] .is_wysiwyg = "true";
defparam \my_reg[30][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N26
cycloneive_lcell_comb \my_reg[18][15]~feeder (
// Equation(s):
// \my_reg[18][15]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat18),
	.cin(gnd),
	.combout(\my_reg[18][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[18][15]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[18][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N27
dffeas \my_reg[18][15] (
	.clk(CLK),
	.d(\my_reg[18][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][15] .is_wysiwyg = "true";
defparam \my_reg[18][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N24
cycloneive_lcell_comb \Mux16~2 (
// Equation(s):
// \Mux16~2_combout  = (dcifimemload_24 & ((\my_reg[26][15]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\my_reg[18][15]~q  & !dcifimemload_23))))

	.dataa(\my_reg[26][15]~q ),
	.datab(\my_reg[18][15]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~2 .lut_mask = 16'hF0AC;
defparam \Mux16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N20
cycloneive_lcell_comb \Mux16~3 (
// Equation(s):
// \Mux16~3_combout  = (dcifimemload_23 & ((\Mux16~2_combout  & ((\my_reg[30][15]~q ))) # (!\Mux16~2_combout  & (\my_reg[22][15]~q )))) # (!dcifimemload_23 & (((\Mux16~2_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[22][15]~q ),
	.datac(\my_reg[30][15]~q ),
	.datad(\Mux16~2_combout ),
	.cin(gnd),
	.combout(\Mux16~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~3 .lut_mask = 16'hF588;
defparam \Mux16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y30_N3
dffeas \my_reg[28][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][15] .is_wysiwyg = "true";
defparam \my_reg[28][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N1
dffeas \my_reg[16][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][15] .is_wysiwyg = "true";
defparam \my_reg[16][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N0
cycloneive_lcell_comb \Mux16~4 (
// Equation(s):
// \Mux16~4_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[24][15]~q )) # (!dcifimemload_24 & ((\my_reg[16][15]~q )))))

	.dataa(\my_reg[24][15]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[16][15]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~4 .lut_mask = 16'hEE30;
defparam \Mux16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N2
cycloneive_lcell_comb \Mux16~5 (
// Equation(s):
// \Mux16~5_combout  = (dcifimemload_23 & ((\Mux16~4_combout  & ((\my_reg[28][15]~q ))) # (!\Mux16~4_combout  & (\my_reg[20][15]~q )))) # (!dcifimemload_23 & (((\Mux16~4_combout ))))

	.dataa(\my_reg[20][15]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[28][15]~q ),
	.datad(\Mux16~4_combout ),
	.cin(gnd),
	.combout(\Mux16~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~5 .lut_mask = 16'hF388;
defparam \Mux16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N26
cycloneive_lcell_comb \Mux16~6 (
// Equation(s):
// \Mux16~6_combout  = (dcifimemload_22 & ((\Mux16~3_combout ) # ((dcifimemload_21)))) # (!dcifimemload_22 & (((!dcifimemload_21 & \Mux16~5_combout ))))

	.dataa(dcifimemload_22),
	.datab(\Mux16~3_combout ),
	.datac(dcifimemload_21),
	.datad(\Mux16~5_combout ),
	.cin(gnd),
	.combout(\Mux16~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~6 .lut_mask = 16'hADA8;
defparam \Mux16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N14
cycloneive_lcell_comb \my_reg[29][15]~feeder (
// Equation(s):
// \my_reg[29][15]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat18),
	.cin(gnd),
	.combout(\my_reg[29][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[29][15]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[29][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N15
dffeas \my_reg[29][15] (
	.clk(CLK),
	.d(\my_reg[29][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][15] .is_wysiwyg = "true";
defparam \my_reg[29][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N29
dffeas \my_reg[17][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][15] .is_wysiwyg = "true";
defparam \my_reg[17][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N28
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (dcifimemload_23 & ((\my_reg[21][15]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[17][15]~q  & !dcifimemload_24))))

	.dataa(\my_reg[21][15]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[17][15]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'hCCB8;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N24
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// \Mux16~1_combout  = (dcifimemload_24 & ((\Mux16~0_combout  & ((\my_reg[29][15]~q ))) # (!\Mux16~0_combout  & (\my_reg[25][15]~q )))) # (!dcifimemload_24 & (((\Mux16~0_combout ))))

	.dataa(\my_reg[25][15]~q ),
	.datab(\my_reg[29][15]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux16~0_combout ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hCFA0;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N8
cycloneive_lcell_comb \Mux16~9 (
// Equation(s):
// \Mux16~9_combout  = (dcifimemload_21 & ((\Mux16~6_combout  & (\Mux16~8_combout )) # (!\Mux16~6_combout  & ((\Mux16~1_combout ))))) # (!dcifimemload_21 & (((\Mux16~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux16~8_combout ),
	.datac(\Mux16~6_combout ),
	.datad(\Mux16~1_combout ),
	.cin(gnd),
	.combout(\Mux16~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~9 .lut_mask = 16'hDAD0;
defparam \Mux16~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N20
cycloneive_lcell_comb \my_reg[15][15]~feeder (
// Equation(s):
// \my_reg[15][15]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat18),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[15][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[15][15]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[15][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N21
dffeas \my_reg[15][15] (
	.clk(CLK),
	.d(\my_reg[15][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][15] .is_wysiwyg = "true";
defparam \my_reg[15][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N6
cycloneive_lcell_comb \my_reg[12][15]~feeder (
// Equation(s):
// \my_reg[12][15]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat18),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[12][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[12][15]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[12][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N7
dffeas \my_reg[12][15] (
	.clk(CLK),
	.d(\my_reg[12][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][15] .is_wysiwyg = "true";
defparam \my_reg[12][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N7
dffeas \my_reg[13][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][15] .is_wysiwyg = "true";
defparam \my_reg[13][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N6
cycloneive_lcell_comb \Mux16~17 (
// Equation(s):
// \Mux16~17_combout  = (dcifimemload_21 & (((\my_reg[13][15]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\my_reg[12][15]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[12][15]~q ),
	.datac(\my_reg[13][15]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux16~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~17 .lut_mask = 16'hAAE4;
defparam \Mux16~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N20
cycloneive_lcell_comb \Mux16~18 (
// Equation(s):
// \Mux16~18_combout  = (\Mux16~17_combout  & (((\my_reg[15][15]~q ) # (!dcifimemload_22)))) # (!\Mux16~17_combout  & (\my_reg[14][15]~q  & ((dcifimemload_22))))

	.dataa(\my_reg[14][15]~q ),
	.datab(\my_reg[15][15]~q ),
	.datac(\Mux16~17_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux16~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~18 .lut_mask = 16'hCAF0;
defparam \Mux16~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N0
cycloneive_lcell_comb \my_reg[9][15]~feeder (
// Equation(s):
// \my_reg[9][15]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat18),
	.cin(gnd),
	.combout(\my_reg[9][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[9][15]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[9][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y31_N1
dffeas \my_reg[9][15] (
	.clk(CLK),
	.d(\my_reg[9][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][15] .is_wysiwyg = "true";
defparam \my_reg[9][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N17
dffeas \my_reg[10][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][15] .is_wysiwyg = "true";
defparam \my_reg[10][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N16
cycloneive_lcell_comb \Mux16~10 (
// Equation(s):
// \Mux16~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[10][15]~q ))) # (!dcifimemload_22 & (\my_reg[8][15]~q ))))

	.dataa(\my_reg[8][15]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[10][15]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux16~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~10 .lut_mask = 16'hFC22;
defparam \Mux16~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N19
dffeas \my_reg[11][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][15] .is_wysiwyg = "true";
defparam \my_reg[11][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N22
cycloneive_lcell_comb \Mux16~11 (
// Equation(s):
// \Mux16~11_combout  = (dcifimemload_21 & ((\Mux16~10_combout  & ((\my_reg[11][15]~q ))) # (!\Mux16~10_combout  & (\my_reg[9][15]~q )))) # (!dcifimemload_21 & (((\Mux16~10_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][15]~q ),
	.datac(\Mux16~10_combout ),
	.datad(\my_reg[11][15]~q ),
	.cin(gnd),
	.combout(\Mux16~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~11 .lut_mask = 16'hF858;
defparam \Mux16~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y37_N9
dffeas \my_reg[3][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][15] .is_wysiwyg = "true";
defparam \my_reg[3][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N8
cycloneive_lcell_comb \Mux16~14 (
// Equation(s):
// \Mux16~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][15]~q ))) # (!dcifimemload_22 & (\my_reg[1][15]~q ))))

	.dataa(\my_reg[1][15]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[3][15]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux16~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~14 .lut_mask = 16'hC088;
defparam \Mux16~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N4
cycloneive_lcell_comb \Mux16~15 (
// Equation(s):
// \Mux16~15_combout  = (\Mux16~14_combout ) # ((\my_reg[2][15]~q  & (dcifimemload_22 & !dcifimemload_21)))

	.dataa(\my_reg[2][15]~q ),
	.datab(dcifimemload_22),
	.datac(dcifimemload_21),
	.datad(\Mux16~14_combout ),
	.cin(gnd),
	.combout(\Mux16~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~15 .lut_mask = 16'hFF08;
defparam \Mux16~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N19
dffeas \my_reg[7][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][15] .is_wysiwyg = "true";
defparam \my_reg[7][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N13
dffeas \my_reg[4][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][15] .is_wysiwyg = "true";
defparam \my_reg[4][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N12
cycloneive_lcell_comb \Mux16~12 (
// Equation(s):
// \Mux16~12_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\my_reg[5][15]~q )) # (!dcifimemload_21 & ((\my_reg[4][15]~q )))))

	.dataa(\my_reg[5][15]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[4][15]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux16~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~12 .lut_mask = 16'hEE30;
defparam \Mux16~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N18
cycloneive_lcell_comb \Mux16~13 (
// Equation(s):
// \Mux16~13_combout  = (dcifimemload_22 & ((\Mux16~12_combout  & ((\my_reg[7][15]~q ))) # (!\Mux16~12_combout  & (\my_reg[6][15]~q )))) # (!dcifimemload_22 & (((\Mux16~12_combout ))))

	.dataa(\my_reg[6][15]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[7][15]~q ),
	.datad(\Mux16~12_combout ),
	.cin(gnd),
	.combout(\Mux16~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~13 .lut_mask = 16'hF388;
defparam \Mux16~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N10
cycloneive_lcell_comb \Mux16~16 (
// Equation(s):
// \Mux16~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & ((\Mux16~13_combout ))) # (!dcifimemload_23 & (\Mux16~15_combout ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux16~15_combout ),
	.datad(\Mux16~13_combout ),
	.cin(gnd),
	.combout(\Mux16~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~16 .lut_mask = 16'hDC98;
defparam \Mux16~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N6
cycloneive_lcell_comb \Mux16~19 (
// Equation(s):
// \Mux16~19_combout  = (dcifimemload_24 & ((\Mux16~16_combout  & (\Mux16~18_combout )) # (!\Mux16~16_combout  & ((\Mux16~11_combout ))))) # (!dcifimemload_24 & (((\Mux16~16_combout ))))

	.dataa(dcifimemload_24),
	.datab(\Mux16~18_combout ),
	.datac(\Mux16~11_combout ),
	.datad(\Mux16~16_combout ),
	.cin(gnd),
	.combout(\Mux16~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~19 .lut_mask = 16'hDDA0;
defparam \Mux16~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y32_N23
dffeas \my_reg[5][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][15] .is_wysiwyg = "true";
defparam \my_reg[5][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N22
cycloneive_lcell_comb \Mux48~0 (
// Equation(s):
// \Mux48~0_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][15]~q ))) # (!dcifimemload_16 & (\my_reg[4][15]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[4][15]~q ),
	.datac(\my_reg[5][15]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux48~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~0 .lut_mask = 16'hFA44;
defparam \Mux48~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y32_N21
dffeas \my_reg[6][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][15] .is_wysiwyg = "true";
defparam \my_reg[6][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N20
cycloneive_lcell_comb \Mux48~1 (
// Equation(s):
// \Mux48~1_combout  = (\Mux48~0_combout  & ((\my_reg[7][15]~q ) # ((!dcifimemload_17)))) # (!\Mux48~0_combout  & (((\my_reg[6][15]~q  & dcifimemload_17))))

	.dataa(\Mux48~0_combout ),
	.datab(\my_reg[7][15]~q ),
	.datac(\my_reg[6][15]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux48~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~1 .lut_mask = 16'hD8AA;
defparam \Mux48~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N20
cycloneive_lcell_comb \my_reg[14][15]~feeder (
// Equation(s):
// \my_reg[14][15]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat18),
	.cin(gnd),
	.combout(\my_reg[14][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[14][15]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[14][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N21
dffeas \my_reg[14][15] (
	.clk(CLK),
	.d(\my_reg[14][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][15] .is_wysiwyg = "true";
defparam \my_reg[14][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N18
cycloneive_lcell_comb \Mux48~7 (
// Equation(s):
// \Mux48~7_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\my_reg[13][15]~q )) # (!dcifimemload_16 & ((\my_reg[12][15]~q )))))

	.dataa(\my_reg[13][15]~q ),
	.datab(\my_reg[12][15]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux48~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~7 .lut_mask = 16'hFA0C;
defparam \Mux48~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N28
cycloneive_lcell_comb \Mux48~8 (
// Equation(s):
// \Mux48~8_combout  = (dcifimemload_17 & ((\Mux48~7_combout  & (\my_reg[15][15]~q )) # (!\Mux48~7_combout  & ((\my_reg[14][15]~q ))))) # (!dcifimemload_17 & (((\Mux48~7_combout ))))

	.dataa(\my_reg[15][15]~q ),
	.datab(\my_reg[14][15]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux48~7_combout ),
	.cin(gnd),
	.combout(\Mux48~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~8 .lut_mask = 16'hAFC0;
defparam \Mux48~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N13
dffeas \my_reg[8][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][15] .is_wysiwyg = "true";
defparam \my_reg[8][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N12
cycloneive_lcell_comb \Mux48~2 (
// Equation(s):
// \Mux48~2_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\my_reg[10][15]~q )) # (!dcifimemload_17 & ((\my_reg[8][15]~q )))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[10][15]~q ),
	.datac(\my_reg[8][15]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux48~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~2 .lut_mask = 16'hEE50;
defparam \Mux48~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N18
cycloneive_lcell_comb \Mux48~3 (
// Equation(s):
// \Mux48~3_combout  = (dcifimemload_16 & ((\Mux48~2_combout  & ((\my_reg[11][15]~q ))) # (!\Mux48~2_combout  & (\my_reg[9][15]~q )))) # (!dcifimemload_16 & (((\Mux48~2_combout ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[9][15]~q ),
	.datac(\my_reg[11][15]~q ),
	.datad(\Mux48~2_combout ),
	.cin(gnd),
	.combout(\Mux48~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~3 .lut_mask = 16'hF588;
defparam \Mux48~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y39_N31
dffeas \my_reg[2][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][15] .is_wysiwyg = "true";
defparam \my_reg[2][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N29
dffeas \my_reg[1][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][15] .is_wysiwyg = "true";
defparam \my_reg[1][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N28
cycloneive_lcell_comb \Mux48~4 (
// Equation(s):
// \Mux48~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\my_reg[3][15]~q )) # (!dcifimemload_17 & ((\my_reg[1][15]~q )))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[3][15]~q ),
	.datac(\my_reg[1][15]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux48~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~4 .lut_mask = 16'hD800;
defparam \Mux48~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N30
cycloneive_lcell_comb \Mux48~5 (
// Equation(s):
// \Mux48~5_combout  = (\Mux48~4_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \my_reg[2][15]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\my_reg[2][15]~q ),
	.datad(\Mux48~4_combout ),
	.cin(gnd),
	.combout(\Mux48~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~5 .lut_mask = 16'hFF20;
defparam \Mux48~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N10
cycloneive_lcell_comb \Mux48~6 (
// Equation(s):
// \Mux48~6_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\Mux48~3_combout )) # (!dcifimemload_19 & ((\Mux48~5_combout )))))

	.dataa(dcifimemload_18),
	.datab(\Mux48~3_combout ),
	.datac(dcifimemload_19),
	.datad(\Mux48~5_combout ),
	.cin(gnd),
	.combout(\Mux48~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~6 .lut_mask = 16'hE5E0;
defparam \Mux48~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N12
cycloneive_lcell_comb \my_reg[23][15]~feeder (
// Equation(s):
// \my_reg[23][15]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat18),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[23][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[23][15]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[23][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N13
dffeas \my_reg[23][15] (
	.clk(CLK),
	.d(\my_reg[23][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][15] .is_wysiwyg = "true";
defparam \my_reg[23][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N18
cycloneive_lcell_comb \Mux48~17 (
// Equation(s):
// \Mux48~17_combout  = (dcifimemload_19 & ((\my_reg[27][15]~q ) # ((dcifimemload_18)))) # (!dcifimemload_19 & (((\my_reg[19][15]~q  & !dcifimemload_18))))

	.dataa(\my_reg[27][15]~q ),
	.datab(\my_reg[19][15]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux48~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~17 .lut_mask = 16'hF0AC;
defparam \Mux48~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N8
cycloneive_lcell_comb \Mux48~18 (
// Equation(s):
// \Mux48~18_combout  = (\Mux48~17_combout  & (((\my_reg[31][15]~q ) # (!dcifimemload_18)))) # (!\Mux48~17_combout  & (\my_reg[23][15]~q  & ((dcifimemload_18))))

	.dataa(\my_reg[23][15]~q ),
	.datab(\Mux48~17_combout ),
	.datac(\my_reg[31][15]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux48~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~18 .lut_mask = 16'hE2CC;
defparam \Mux48~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N12
cycloneive_lcell_comb \my_reg[24][15]~feeder (
// Equation(s):
// \my_reg[24][15]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat18),
	.cin(gnd),
	.combout(\my_reg[24][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[24][15]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[24][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y30_N13
dffeas \my_reg[24][15] (
	.clk(CLK),
	.d(\my_reg[24][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][15] .is_wysiwyg = "true";
defparam \my_reg[24][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N8
cycloneive_lcell_comb \Mux48~15 (
// Equation(s):
// \Mux48~15_combout  = (\Mux48~14_combout  & (((\my_reg[28][15]~q ) # (!dcifimemload_19)))) # (!\Mux48~14_combout  & (\my_reg[24][15]~q  & (dcifimemload_19)))

	.dataa(\Mux48~14_combout ),
	.datab(\my_reg[24][15]~q ),
	.datac(dcifimemload_19),
	.datad(\my_reg[28][15]~q ),
	.cin(gnd),
	.combout(\Mux48~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~15 .lut_mask = 16'hEA4A;
defparam \Mux48~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N31
dffeas \my_reg[26][15] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][15] .is_wysiwyg = "true";
defparam \my_reg[26][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N20
cycloneive_lcell_comb \Mux48~12 (
// Equation(s):
// \Mux48~12_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[22][15]~q ))) # (!dcifimemload_18 & (\my_reg[18][15]~q ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[18][15]~q ),
	.datac(\my_reg[22][15]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux48~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~12 .lut_mask = 16'hFA44;
defparam \Mux48~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N30
cycloneive_lcell_comb \Mux48~13 (
// Equation(s):
// \Mux48~13_combout  = (dcifimemload_19 & ((\Mux48~12_combout  & (\my_reg[30][15]~q )) # (!\Mux48~12_combout  & ((\my_reg[26][15]~q ))))) # (!dcifimemload_19 & (((\Mux48~12_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[30][15]~q ),
	.datac(\my_reg[26][15]~q ),
	.datad(\Mux48~12_combout ),
	.cin(gnd),
	.combout(\Mux48~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~13 .lut_mask = 16'hDDA0;
defparam \Mux48~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N14
cycloneive_lcell_comb \Mux48~16 (
// Equation(s):
// \Mux48~16_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux48~13_combout ))) # (!dcifimemload_17 & (\Mux48~15_combout ))))

	.dataa(dcifimemload_16),
	.datab(\Mux48~15_combout ),
	.datac(dcifimemload_17),
	.datad(\Mux48~13_combout ),
	.cin(gnd),
	.combout(\Mux48~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~16 .lut_mask = 16'hF4A4;
defparam \Mux48~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N10
cycloneive_lcell_comb \my_reg[21][15]~feeder (
// Equation(s):
// \my_reg[21][15]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat18),
	.cin(gnd),
	.combout(\my_reg[21][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][15]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[21][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N11
dffeas \my_reg[21][15] (
	.clk(CLK),
	.d(\my_reg[21][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][15] .is_wysiwyg = "true";
defparam \my_reg[21][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N24
cycloneive_lcell_comb \my_reg[25][15]~feeder (
// Equation(s):
// \my_reg[25][15]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat18),
	.cin(gnd),
	.combout(\my_reg[25][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][15]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[25][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N25
dffeas \my_reg[25][15] (
	.clk(CLK),
	.d(\my_reg[25][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][15] .is_wysiwyg = "true";
defparam \my_reg[25][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N20
cycloneive_lcell_comb \Mux48~10 (
// Equation(s):
// \Mux48~10_combout  = (dcifimemload_19 & (((\my_reg[25][15]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[17][15]~q  & ((!dcifimemload_18))))

	.dataa(\my_reg[17][15]~q ),
	.datab(\my_reg[25][15]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux48~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~10 .lut_mask = 16'hF0CA;
defparam \Mux48~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N26
cycloneive_lcell_comb \Mux48~11 (
// Equation(s):
// \Mux48~11_combout  = (dcifimemload_18 & ((\Mux48~10_combout  & ((\my_reg[29][15]~q ))) # (!\Mux48~10_combout  & (\my_reg[21][15]~q )))) # (!dcifimemload_18 & (((\Mux48~10_combout ))))

	.dataa(\my_reg[21][15]~q ),
	.datab(\my_reg[29][15]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux48~10_combout ),
	.cin(gnd),
	.combout(\Mux48~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~11 .lut_mask = 16'hCFA0;
defparam \Mux48~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N28
cycloneive_lcell_comb \my_reg[14][14]~feeder (
// Equation(s):
// \my_reg[14][14]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat19),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[14][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[14][14]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[14][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N29
dffeas \my_reg[14][14] (
	.clk(CLK),
	.d(\my_reg[14][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][14] .is_wysiwyg = "true";
defparam \my_reg[14][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N29
dffeas \my_reg[12][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][14] .is_wysiwyg = "true";
defparam \my_reg[12][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N13
dffeas \my_reg[13][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][14] .is_wysiwyg = "true";
defparam \my_reg[13][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N12
cycloneive_lcell_comb \Mux17~17 (
// Equation(s):
// \Mux17~17_combout  = (dcifimemload_21 & (((\my_reg[13][14]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\my_reg[12][14]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[12][14]~q ),
	.datac(\my_reg[13][14]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux17~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~17 .lut_mask = 16'hAAE4;
defparam \Mux17~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N26
cycloneive_lcell_comb \Mux17~18 (
// Equation(s):
// \Mux17~18_combout  = (dcifimemload_22 & ((\Mux17~17_combout  & (\my_reg[15][14]~q )) # (!\Mux17~17_combout  & ((\my_reg[14][14]~q ))))) # (!dcifimemload_22 & (((\Mux17~17_combout ))))

	.dataa(\my_reg[15][14]~q ),
	.datab(\my_reg[14][14]~q ),
	.datac(dcifimemload_22),
	.datad(\Mux17~17_combout ),
	.cin(gnd),
	.combout(\Mux17~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~18 .lut_mask = 16'hAFC0;
defparam \Mux17~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N22
cycloneive_lcell_comb \my_reg[7][14]~feeder (
// Equation(s):
// \my_reg[7][14]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat19),
	.cin(gnd),
	.combout(\my_reg[7][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[7][14]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[7][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y43_N23
dffeas \my_reg[7][14] (
	.clk(CLK),
	.d(\my_reg[7][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][14] .is_wysiwyg = "true";
defparam \my_reg[7][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N5
dffeas \my_reg[4][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][14] .is_wysiwyg = "true";
defparam \my_reg[4][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N22
cycloneive_lcell_comb \Mux17~10 (
// Equation(s):
// \Mux17~10_combout  = (dcifimemload_21 & ((\my_reg[5][14]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[4][14]~q  & !dcifimemload_22))))

	.dataa(\my_reg[5][14]~q ),
	.datab(\my_reg[4][14]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux17~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~10 .lut_mask = 16'hF0AC;
defparam \Mux17~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N28
cycloneive_lcell_comb \Mux17~11 (
// Equation(s):
// \Mux17~11_combout  = (\Mux17~10_combout  & (((\my_reg[7][14]~q ) # (!dcifimemload_22)))) # (!\Mux17~10_combout  & (\my_reg[6][14]~q  & ((dcifimemload_22))))

	.dataa(\my_reg[6][14]~q ),
	.datab(\my_reg[7][14]~q ),
	.datac(\Mux17~10_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux17~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~11 .lut_mask = 16'hCAF0;
defparam \Mux17~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y40_N1
dffeas \my_reg[2][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][14] .is_wysiwyg = "true";
defparam \my_reg[2][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y40_N3
dffeas \my_reg[1][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][14] .is_wysiwyg = "true";
defparam \my_reg[1][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y42_N31
dffeas \my_reg[3][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][14] .is_wysiwyg = "true";
defparam \my_reg[3][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N30
cycloneive_lcell_comb \Mux17~14 (
// Equation(s):
// \Mux17~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][14]~q ))) # (!dcifimemload_22 & (\my_reg[1][14]~q ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[1][14]~q ),
	.datac(\my_reg[3][14]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux17~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~14 .lut_mask = 16'hA088;
defparam \Mux17~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N30
cycloneive_lcell_comb \Mux17~15 (
// Equation(s):
// \Mux17~15_combout  = (\Mux17~14_combout ) # ((dcifimemload_22 & (\my_reg[2][14]~q  & !dcifimemload_21)))

	.dataa(dcifimemload_22),
	.datab(\my_reg[2][14]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux17~14_combout ),
	.cin(gnd),
	.combout(\Mux17~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~15 .lut_mask = 16'hFF08;
defparam \Mux17~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y30_N15
dffeas \my_reg[9][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][14] .is_wysiwyg = "true";
defparam \my_reg[9][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N25
dffeas \my_reg[11][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][14] .is_wysiwyg = "true";
defparam \my_reg[11][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N7
dffeas \my_reg[8][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][14] .is_wysiwyg = "true";
defparam \my_reg[8][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N6
cycloneive_lcell_comb \Mux17~12 (
// Equation(s):
// \Mux17~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][14]~q )) # (!dcifimemload_22 & ((\my_reg[8][14]~q )))))

	.dataa(\my_reg[10][14]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[8][14]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux17~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~12 .lut_mask = 16'hEE30;
defparam \Mux17~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N24
cycloneive_lcell_comb \Mux17~13 (
// Equation(s):
// \Mux17~13_combout  = (dcifimemload_21 & ((\Mux17~12_combout  & ((\my_reg[11][14]~q ))) # (!\Mux17~12_combout  & (\my_reg[9][14]~q )))) # (!dcifimemload_21 & (((\Mux17~12_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][14]~q ),
	.datac(\my_reg[11][14]~q ),
	.datad(\Mux17~12_combout ),
	.cin(gnd),
	.combout(\Mux17~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~13 .lut_mask = 16'hF588;
defparam \Mux17~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N12
cycloneive_lcell_comb \Mux17~16 (
// Equation(s):
// \Mux17~16_combout  = (dcifimemload_23 & (dcifimemload_24)) # (!dcifimemload_23 & ((dcifimemload_24 & ((\Mux17~13_combout ))) # (!dcifimemload_24 & (\Mux17~15_combout ))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux17~15_combout ),
	.datad(\Mux17~13_combout ),
	.cin(gnd),
	.combout(\Mux17~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~16 .lut_mask = 16'hDC98;
defparam \Mux17~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N8
cycloneive_lcell_comb \Mux17~19 (
// Equation(s):
// \Mux17~19_combout  = (dcifimemload_23 & ((\Mux17~16_combout  & (\Mux17~18_combout )) # (!\Mux17~16_combout  & ((\Mux17~11_combout ))))) # (!dcifimemload_23 & (((\Mux17~16_combout ))))

	.dataa(\Mux17~18_combout ),
	.datab(dcifimemload_23),
	.datac(\Mux17~11_combout ),
	.datad(\Mux17~16_combout ),
	.cin(gnd),
	.combout(\Mux17~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~19 .lut_mask = 16'hBBC0;
defparam \Mux17~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N29
dffeas \my_reg[21][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][14] .is_wysiwyg = "true";
defparam \my_reg[21][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N9
dffeas \my_reg[29][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][14] .is_wysiwyg = "true";
defparam \my_reg[29][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N8
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// \Mux17~1_combout  = (\Mux17~0_combout  & (((\my_reg[29][14]~q ) # (!dcifimemload_23)))) # (!\Mux17~0_combout  & (\my_reg[21][14]~q  & ((dcifimemload_23))))

	.dataa(\Mux17~0_combout ),
	.datab(\my_reg[21][14]~q ),
	.datac(\my_reg[29][14]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hE4AA;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N28
cycloneive_lcell_comb \my_reg[31][14]~feeder (
// Equation(s):
// \my_reg[31][14]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat19),
	.cin(gnd),
	.combout(\my_reg[31][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[31][14]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[31][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N29
dffeas \my_reg[31][14] (
	.clk(CLK),
	.d(\my_reg[31][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][14] .is_wysiwyg = "true";
defparam \my_reg[31][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N9
dffeas \my_reg[27][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][14] .is_wysiwyg = "true";
defparam \my_reg[27][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N4
cycloneive_lcell_comb \Mux17~7 (
// Equation(s):
// \Mux17~7_combout  = (dcifimemload_24 & (((\my_reg[27][14]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\my_reg[19][14]~q  & ((!dcifimemload_23))))

	.dataa(\my_reg[19][14]~q ),
	.datab(\my_reg[27][14]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux17~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~7 .lut_mask = 16'hF0CA;
defparam \Mux17~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N26
cycloneive_lcell_comb \Mux17~8 (
// Equation(s):
// \Mux17~8_combout  = (dcifimemload_23 & ((\Mux17~7_combout  & ((\my_reg[31][14]~q ))) # (!\Mux17~7_combout  & (\my_reg[23][14]~q )))) # (!dcifimemload_23 & (((\Mux17~7_combout ))))

	.dataa(\my_reg[23][14]~q ),
	.datab(\my_reg[31][14]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux17~7_combout ),
	.cin(gnd),
	.combout(\Mux17~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~8 .lut_mask = 16'hCFA0;
defparam \Mux17~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y30_N19
dffeas \my_reg[28][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][14] .is_wysiwyg = "true";
defparam \my_reg[28][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N13
dffeas \my_reg[16][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][14] .is_wysiwyg = "true";
defparam \my_reg[16][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N12
cycloneive_lcell_comb \Mux17~4 (
// Equation(s):
// \Mux17~4_combout  = (dcifimemload_23 & ((\my_reg[20][14]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[16][14]~q  & !dcifimemload_24))))

	.dataa(\my_reg[20][14]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[16][14]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~4 .lut_mask = 16'hCCB8;
defparam \Mux17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N18
cycloneive_lcell_comb \Mux17~5 (
// Equation(s):
// \Mux17~5_combout  = (dcifimemload_24 & ((\Mux17~4_combout  & ((\my_reg[28][14]~q ))) # (!\Mux17~4_combout  & (\my_reg[24][14]~q )))) # (!dcifimemload_24 & (((\Mux17~4_combout ))))

	.dataa(\my_reg[24][14]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[28][14]~q ),
	.datad(\Mux17~4_combout ),
	.cin(gnd),
	.combout(\Mux17~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~5 .lut_mask = 16'hF388;
defparam \Mux17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y30_N11
dffeas \my_reg[26][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][14] .is_wysiwyg = "true";
defparam \my_reg[26][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N18
cycloneive_lcell_comb \my_reg[30][14]~feeder (
// Equation(s):
// \my_reg[30][14]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat19),
	.cin(gnd),
	.combout(\my_reg[30][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[30][14]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[30][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N19
dffeas \my_reg[30][14] (
	.clk(CLK),
	.d(\my_reg[30][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][14] .is_wysiwyg = "true";
defparam \my_reg[30][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N13
dffeas \my_reg[18][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][14] .is_wysiwyg = "true";
defparam \my_reg[18][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N12
cycloneive_lcell_comb \Mux17~2 (
// Equation(s):
// \Mux17~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[22][14]~q )) # (!dcifimemload_23 & ((\my_reg[18][14]~q )))))

	.dataa(\my_reg[22][14]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[18][14]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~2 .lut_mask = 16'hEE30;
defparam \Mux17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N0
cycloneive_lcell_comb \Mux17~3 (
// Equation(s):
// \Mux17~3_combout  = (dcifimemload_24 & ((\Mux17~2_combout  & ((\my_reg[30][14]~q ))) # (!\Mux17~2_combout  & (\my_reg[26][14]~q )))) # (!dcifimemload_24 & (((\Mux17~2_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[26][14]~q ),
	.datac(\my_reg[30][14]~q ),
	.datad(\Mux17~2_combout ),
	.cin(gnd),
	.combout(\Mux17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~3 .lut_mask = 16'hF588;
defparam \Mux17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N18
cycloneive_lcell_comb \Mux17~6 (
// Equation(s):
// \Mux17~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux17~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & (\Mux17~5_combout )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux17~5_combout ),
	.datad(\Mux17~3_combout ),
	.cin(gnd),
	.combout(\Mux17~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~6 .lut_mask = 16'hBA98;
defparam \Mux17~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N28
cycloneive_lcell_comb \Mux17~9 (
// Equation(s):
// \Mux17~9_combout  = (dcifimemload_21 & ((\Mux17~6_combout  & ((\Mux17~8_combout ))) # (!\Mux17~6_combout  & (\Mux17~1_combout )))) # (!dcifimemload_21 & (((\Mux17~6_combout ))))

	.dataa(\Mux17~1_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux17~8_combout ),
	.datad(\Mux17~6_combout ),
	.cin(gnd),
	.combout(\Mux17~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~9 .lut_mask = 16'hF388;
defparam \Mux17~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N26
cycloneive_lcell_comb \my_reg[15][14]~feeder (
// Equation(s):
// \my_reg[15][14]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat19),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[15][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[15][14]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[15][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N27
dffeas \my_reg[15][14] (
	.clk(CLK),
	.d(\my_reg[15][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][14] .is_wysiwyg = "true";
defparam \my_reg[15][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N28
cycloneive_lcell_comb \Mux49~7 (
// Equation(s):
// \Mux49~7_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\my_reg[13][14]~q )) # (!dcifimemload_16 & ((\my_reg[12][14]~q )))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[13][14]~q ),
	.datac(\my_reg[12][14]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux49~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~7 .lut_mask = 16'hEE50;
defparam \Mux49~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N2
cycloneive_lcell_comb \Mux49~8 (
// Equation(s):
// \Mux49~8_combout  = (dcifimemload_17 & ((\Mux49~7_combout  & (\my_reg[15][14]~q )) # (!\Mux49~7_combout  & ((\my_reg[14][14]~q ))))) # (!dcifimemload_17 & (((\Mux49~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[15][14]~q ),
	.datac(\my_reg[14][14]~q ),
	.datad(\Mux49~7_combout ),
	.cin(gnd),
	.combout(\Mux49~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~8 .lut_mask = 16'hDDA0;
defparam \Mux49~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y30_N29
dffeas \my_reg[10][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][14] .is_wysiwyg = "true";
defparam \my_reg[10][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N28
cycloneive_lcell_comb \Mux49~0 (
// Equation(s):
// \Mux49~0_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[10][14]~q ))) # (!dcifimemload_17 & (\my_reg[8][14]~q ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[8][14]~q ),
	.datac(\my_reg[10][14]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux49~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~0 .lut_mask = 16'hFA44;
defparam \Mux49~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N14
cycloneive_lcell_comb \Mux49~1 (
// Equation(s):
// \Mux49~1_combout  = (dcifimemload_16 & ((\Mux49~0_combout  & (\my_reg[11][14]~q )) # (!\Mux49~0_combout  & ((\my_reg[9][14]~q ))))) # (!dcifimemload_16 & (((\Mux49~0_combout ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[11][14]~q ),
	.datac(\my_reg[9][14]~q ),
	.datad(\Mux49~0_combout ),
	.cin(gnd),
	.combout(\Mux49~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~1 .lut_mask = 16'hDDA0;
defparam \Mux49~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N12
cycloneive_lcell_comb \my_reg[6][14]~feeder (
// Equation(s):
// \my_reg[6][14]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat19),
	.cin(gnd),
	.combout(\my_reg[6][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[6][14]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[6][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y43_N13
dffeas \my_reg[6][14] (
	.clk(CLK),
	.d(\my_reg[6][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][14] .is_wysiwyg = "true";
defparam \my_reg[6][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N4
cycloneive_lcell_comb \Mux49~2 (
// Equation(s):
// \Mux49~2_combout  = (dcifimemload_16 & ((\my_reg[5][14]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\my_reg[4][14]~q  & !dcifimemload_17))))

	.dataa(\my_reg[5][14]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[4][14]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux49~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~2 .lut_mask = 16'hCCB8;
defparam \Mux49~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N26
cycloneive_lcell_comb \Mux49~3 (
// Equation(s):
// \Mux49~3_combout  = (\Mux49~2_combout  & ((\my_reg[7][14]~q ) # ((!dcifimemload_17)))) # (!\Mux49~2_combout  & (((\my_reg[6][14]~q  & dcifimemload_17))))

	.dataa(\my_reg[7][14]~q ),
	.datab(\my_reg[6][14]~q ),
	.datac(\Mux49~2_combout ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux49~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~3 .lut_mask = 16'hACF0;
defparam \Mux49~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N2
cycloneive_lcell_comb \Mux49~4 (
// Equation(s):
// \Mux49~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\my_reg[3][14]~q )) # (!dcifimemload_17 & ((\my_reg[1][14]~q )))))

	.dataa(\my_reg[3][14]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[1][14]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux49~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~4 .lut_mask = 16'h88C0;
defparam \Mux49~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N0
cycloneive_lcell_comb \Mux49~5 (
// Equation(s):
// \Mux49~5_combout  = (\Mux49~4_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \my_reg[2][14]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\my_reg[2][14]~q ),
	.datad(\Mux49~4_combout ),
	.cin(gnd),
	.combout(\Mux49~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~5 .lut_mask = 16'hFF20;
defparam \Mux49~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N2
cycloneive_lcell_comb \Mux49~6 (
// Equation(s):
// \Mux49~6_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & (\Mux49~3_combout )) # (!dcifimemload_18 & ((\Mux49~5_combout )))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux49~3_combout ),
	.datad(\Mux49~5_combout ),
	.cin(gnd),
	.combout(\Mux49~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~6 .lut_mask = 16'hD9C8;
defparam \Mux49~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N8
cycloneive_lcell_comb \my_reg[25][14]~feeder (
// Equation(s):
// \my_reg[25][14]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat19),
	.cin(gnd),
	.combout(\my_reg[25][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][14]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[25][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N9
dffeas \my_reg[25][14] (
	.clk(CLK),
	.d(\my_reg[25][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][14] .is_wysiwyg = "true";
defparam \my_reg[25][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N28
cycloneive_lcell_comb \Mux49~10 (
// Equation(s):
// \Mux49~10_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[21][14]~q ))) # (!dcifimemload_18 & (\my_reg[17][14]~q ))))

	.dataa(\my_reg[17][14]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[21][14]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux49~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~10 .lut_mask = 16'hFC22;
defparam \Mux49~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N26
cycloneive_lcell_comb \Mux49~11 (
// Equation(s):
// \Mux49~11_combout  = (dcifimemload_19 & ((\Mux49~10_combout  & (\my_reg[29][14]~q )) # (!\Mux49~10_combout  & ((\my_reg[25][14]~q ))))) # (!dcifimemload_19 & (((\Mux49~10_combout ))))

	.dataa(\my_reg[29][14]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[25][14]~q ),
	.datad(\Mux49~10_combout ),
	.cin(gnd),
	.combout(\Mux49~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~11 .lut_mask = 16'hBBC0;
defparam \Mux49~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y30_N21
dffeas \my_reg[20][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][14] .is_wysiwyg = "true";
defparam \my_reg[20][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N20
cycloneive_lcell_comb \Mux49~15 (
// Equation(s):
// \Mux49~15_combout  = (\Mux49~14_combout  & (((\my_reg[28][14]~q )) # (!dcifimemload_18))) # (!\Mux49~14_combout  & (dcifimemload_18 & (\my_reg[20][14]~q )))

	.dataa(\Mux49~14_combout ),
	.datab(dcifimemload_18),
	.datac(\my_reg[20][14]~q ),
	.datad(\my_reg[28][14]~q ),
	.cin(gnd),
	.combout(\Mux49~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~15 .lut_mask = 16'hEA62;
defparam \Mux49~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N10
cycloneive_lcell_comb \Mux49~12 (
// Equation(s):
// \Mux49~12_combout  = (dcifimemload_19 & (((\my_reg[26][14]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[18][14]~q  & ((!dcifimemload_18))))

	.dataa(\my_reg[18][14]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[26][14]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux49~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~12 .lut_mask = 16'hCCE2;
defparam \Mux49~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N27
dffeas \my_reg[22][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][14] .is_wysiwyg = "true";
defparam \my_reg[22][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N28
cycloneive_lcell_comb \Mux49~13 (
// Equation(s):
// \Mux49~13_combout  = (dcifimemload_18 & ((\Mux49~12_combout  & (\my_reg[30][14]~q )) # (!\Mux49~12_combout  & ((\my_reg[22][14]~q ))))) # (!dcifimemload_18 & (((\Mux49~12_combout ))))

	.dataa(\my_reg[30][14]~q ),
	.datab(dcifimemload_18),
	.datac(\Mux49~12_combout ),
	.datad(\my_reg[22][14]~q ),
	.cin(gnd),
	.combout(\Mux49~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~13 .lut_mask = 16'hBCB0;
defparam \Mux49~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N26
cycloneive_lcell_comb \Mux49~16 (
// Equation(s):
// \Mux49~16_combout  = (dcifimemload_17 & (((dcifimemload_16) # (\Mux49~13_combout )))) # (!dcifimemload_17 & (\Mux49~15_combout  & (!dcifimemload_16)))

	.dataa(dcifimemload_17),
	.datab(\Mux49~15_combout ),
	.datac(dcifimemload_16),
	.datad(\Mux49~13_combout ),
	.cin(gnd),
	.combout(\Mux49~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~16 .lut_mask = 16'hAEA4;
defparam \Mux49~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N22
cycloneive_lcell_comb \my_reg[19][14]~feeder (
// Equation(s):
// \my_reg[19][14]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat19),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[19][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[19][14]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[19][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y34_N23
dffeas \my_reg[19][14] (
	.clk(CLK),
	.d(\my_reg[19][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][14] .is_wysiwyg = "true";
defparam \my_reg[19][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N5
dffeas \my_reg[23][14] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][14] .is_wysiwyg = "true";
defparam \my_reg[23][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N4
cycloneive_lcell_comb \Mux49~17 (
// Equation(s):
// \Mux49~17_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[23][14]~q ))) # (!dcifimemload_18 & (\my_reg[19][14]~q ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[19][14]~q ),
	.datac(\my_reg[23][14]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux49~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~17 .lut_mask = 16'hFA44;
defparam \Mux49~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N8
cycloneive_lcell_comb \Mux49~18 (
// Equation(s):
// \Mux49~18_combout  = (dcifimemload_19 & ((\Mux49~17_combout  & (\my_reg[31][14]~q )) # (!\Mux49~17_combout  & ((\my_reg[27][14]~q ))))) # (!dcifimemload_19 & (((\Mux49~17_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[31][14]~q ),
	.datac(\my_reg[27][14]~q ),
	.datad(\Mux49~17_combout ),
	.cin(gnd),
	.combout(\Mux49~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~18 .lut_mask = 16'hDDA0;
defparam \Mux49~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N28
cycloneive_lcell_comb \my_reg[9][13]~feeder (
// Equation(s):
// \my_reg[9][13]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat20),
	.cin(gnd),
	.combout(\my_reg[9][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[9][13]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[9][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N29
dffeas \my_reg[9][13] (
	.clk(CLK),
	.d(\my_reg[9][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][13] .is_wysiwyg = "true";
defparam \my_reg[9][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N25
dffeas \my_reg[8][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][13] .is_wysiwyg = "true";
defparam \my_reg[8][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N8
cycloneive_lcell_comb \Mux18~10 (
// Equation(s):
// \Mux18~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][13]~q )) # (!dcifimemload_22 & ((\my_reg[8][13]~q )))))

	.dataa(\my_reg[10][13]~q ),
	.datab(\my_reg[8][13]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux18~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~10 .lut_mask = 16'hFA0C;
defparam \Mux18~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N10
cycloneive_lcell_comb \Mux18~11 (
// Equation(s):
// \Mux18~11_combout  = (dcifimemload_21 & ((\Mux18~10_combout  & (\my_reg[11][13]~q )) # (!\Mux18~10_combout  & ((\my_reg[9][13]~q ))))) # (!dcifimemload_21 & (((\Mux18~10_combout ))))

	.dataa(\my_reg[11][13]~q ),
	.datab(\my_reg[9][13]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux18~10_combout ),
	.cin(gnd),
	.combout(\Mux18~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~11 .lut_mask = 16'hAFC0;
defparam \Mux18~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N17
dffeas \my_reg[2][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][13] .is_wysiwyg = "true";
defparam \my_reg[2][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N30
cycloneive_lcell_comb \Mux18~15 (
// Equation(s):
// \Mux18~15_combout  = (\Mux18~14_combout ) # ((\my_reg[2][13]~q  & (dcifimemload_22 & !dcifimemload_21)))

	.dataa(\Mux18~14_combout ),
	.datab(\my_reg[2][13]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux18~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~15 .lut_mask = 16'hAAEA;
defparam \Mux18~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y32_N5
dffeas \my_reg[6][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][13] .is_wysiwyg = "true";
defparam \my_reg[6][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N7
dffeas \my_reg[7][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][13] .is_wysiwyg = "true";
defparam \my_reg[7][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N21
dffeas \my_reg[4][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][13] .is_wysiwyg = "true";
defparam \my_reg[4][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N20
cycloneive_lcell_comb \Mux18~12 (
// Equation(s):
// \Mux18~12_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\my_reg[5][13]~q )) # (!dcifimemload_21 & ((\my_reg[4][13]~q )))))

	.dataa(\my_reg[5][13]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[4][13]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux18~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~12 .lut_mask = 16'hEE30;
defparam \Mux18~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N6
cycloneive_lcell_comb \Mux18~13 (
// Equation(s):
// \Mux18~13_combout  = (dcifimemload_22 & ((\Mux18~12_combout  & ((\my_reg[7][13]~q ))) # (!\Mux18~12_combout  & (\my_reg[6][13]~q )))) # (!dcifimemload_22 & (((\Mux18~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[6][13]~q ),
	.datac(\my_reg[7][13]~q ),
	.datad(\Mux18~12_combout ),
	.cin(gnd),
	.combout(\Mux18~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~13 .lut_mask = 16'hF588;
defparam \Mux18~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N8
cycloneive_lcell_comb \Mux18~16 (
// Equation(s):
// \Mux18~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & ((\Mux18~13_combout ))) # (!dcifimemload_23 & (\Mux18~15_combout ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux18~15_combout ),
	.datad(\Mux18~13_combout ),
	.cin(gnd),
	.combout(\Mux18~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~16 .lut_mask = 16'hDC98;
defparam \Mux18~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N9
dffeas \my_reg[14][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][13] .is_wysiwyg = "true";
defparam \my_reg[14][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N18
cycloneive_lcell_comb \my_reg[13][13]~feeder (
// Equation(s):
// \my_reg[13][13]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat20),
	.cin(gnd),
	.combout(\my_reg[13][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[13][13]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[13][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N19
dffeas \my_reg[13][13] (
	.clk(CLK),
	.d(\my_reg[13][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][13] .is_wysiwyg = "true";
defparam \my_reg[13][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N4
cycloneive_lcell_comb \Mux18~17 (
// Equation(s):
// \Mux18~17_combout  = (dcifimemload_21 & (((\my_reg[13][13]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\my_reg[12][13]~q  & ((!dcifimemload_22))))

	.dataa(\my_reg[12][13]~q ),
	.datab(\my_reg[13][13]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux18~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~17 .lut_mask = 16'hF0CA;
defparam \Mux18~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N8
cycloneive_lcell_comb \Mux18~18 (
// Equation(s):
// \Mux18~18_combout  = (dcifimemload_22 & ((\Mux18~17_combout  & (\my_reg[15][13]~q )) # (!\Mux18~17_combout  & ((\my_reg[14][13]~q ))))) # (!dcifimemload_22 & (((\Mux18~17_combout ))))

	.dataa(\my_reg[15][13]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[14][13]~q ),
	.datad(\Mux18~17_combout ),
	.cin(gnd),
	.combout(\Mux18~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~18 .lut_mask = 16'hBBC0;
defparam \Mux18~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N26
cycloneive_lcell_comb \Mux18~19 (
// Equation(s):
// \Mux18~19_combout  = (dcifimemload_24 & ((\Mux18~16_combout  & ((\Mux18~18_combout ))) # (!\Mux18~16_combout  & (\Mux18~11_combout )))) # (!dcifimemload_24 & (((\Mux18~16_combout ))))

	.dataa(dcifimemload_24),
	.datab(\Mux18~11_combout ),
	.datac(\Mux18~16_combout ),
	.datad(\Mux18~18_combout ),
	.cin(gnd),
	.combout(\Mux18~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~19 .lut_mask = 16'hF858;
defparam \Mux18~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N19
dffeas \my_reg[16][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][13] .is_wysiwyg = "true";
defparam \my_reg[16][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N18
cycloneive_lcell_comb \Mux18~4 (
// Equation(s):
// \Mux18~4_combout  = (dcifimemload_24 & ((\my_reg[24][13]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\my_reg[16][13]~q  & !dcifimemload_23))))

	.dataa(\my_reg[24][13]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[16][13]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~4 .lut_mask = 16'hCCB8;
defparam \Mux18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N25
dffeas \my_reg[20][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][13] .is_wysiwyg = "true";
defparam \my_reg[20][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N0
cycloneive_lcell_comb \Mux18~5 (
// Equation(s):
// \Mux18~5_combout  = (\Mux18~4_combout  & ((\my_reg[28][13]~q ) # ((!dcifimemload_23)))) # (!\Mux18~4_combout  & (((\my_reg[20][13]~q  & dcifimemload_23))))

	.dataa(\my_reg[28][13]~q ),
	.datab(\Mux18~4_combout ),
	.datac(\my_reg[20][13]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux18~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~5 .lut_mask = 16'hB8CC;
defparam \Mux18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N22
cycloneive_lcell_comb \Mux18~6 (
// Equation(s):
// \Mux18~6_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\Mux18~3_combout )) # (!dcifimemload_22 & ((\Mux18~5_combout )))))

	.dataa(\Mux18~3_combout ),
	.datab(dcifimemload_21),
	.datac(dcifimemload_22),
	.datad(\Mux18~5_combout ),
	.cin(gnd),
	.combout(\Mux18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~6 .lut_mask = 16'hE3E0;
defparam \Mux18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N1
dffeas \my_reg[29][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][13] .is_wysiwyg = "true";
defparam \my_reg[29][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N26
cycloneive_lcell_comb \my_reg[17][13]~feeder (
// Equation(s):
// \my_reg[17][13]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat20),
	.cin(gnd),
	.combout(\my_reg[17][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[17][13]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[17][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N27
dffeas \my_reg[17][13] (
	.clk(CLK),
	.d(\my_reg[17][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][13] .is_wysiwyg = "true";
defparam \my_reg[17][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N8
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (dcifimemload_23 & ((\my_reg[21][13]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[17][13]~q  & !dcifimemload_24))))

	.dataa(\my_reg[21][13]~q ),
	.datab(\my_reg[17][13]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hF0AC;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N0
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// \Mux18~1_combout  = (dcifimemload_24 & ((\Mux18~0_combout  & ((\my_reg[29][13]~q ))) # (!\Mux18~0_combout  & (\my_reg[25][13]~q )))) # (!dcifimemload_24 & (((\Mux18~0_combout ))))

	.dataa(\my_reg[25][13]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[29][13]~q ),
	.datad(\Mux18~0_combout ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'hF388;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N1
dffeas \my_reg[27][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][13] .is_wysiwyg = "true";
defparam \my_reg[27][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N9
dffeas \my_reg[31][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][13] .is_wysiwyg = "true";
defparam \my_reg[31][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N14
cycloneive_lcell_comb \my_reg[19][13]~feeder (
// Equation(s):
// \my_reg[19][13]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat20),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[19][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[19][13]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[19][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N15
dffeas \my_reg[19][13] (
	.clk(CLK),
	.d(\my_reg[19][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][13] .is_wysiwyg = "true";
defparam \my_reg[19][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N8
cycloneive_lcell_comb \Mux18~7 (
// Equation(s):
// \Mux18~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[23][13]~q )) # (!dcifimemload_23 & ((\my_reg[19][13]~q )))))

	.dataa(\my_reg[23][13]~q ),
	.datab(\my_reg[19][13]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux18~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~7 .lut_mask = 16'hFA0C;
defparam \Mux18~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N8
cycloneive_lcell_comb \Mux18~8 (
// Equation(s):
// \Mux18~8_combout  = (dcifimemload_24 & ((\Mux18~7_combout  & ((\my_reg[31][13]~q ))) # (!\Mux18~7_combout  & (\my_reg[27][13]~q )))) # (!dcifimemload_24 & (((\Mux18~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[27][13]~q ),
	.datac(\my_reg[31][13]~q ),
	.datad(\Mux18~7_combout ),
	.cin(gnd),
	.combout(\Mux18~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~8 .lut_mask = 16'hF588;
defparam \Mux18~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N24
cycloneive_lcell_comb \Mux18~9 (
// Equation(s):
// \Mux18~9_combout  = (\Mux18~6_combout  & (((\Mux18~8_combout )) # (!dcifimemload_21))) # (!\Mux18~6_combout  & (dcifimemload_21 & (\Mux18~1_combout )))

	.dataa(\Mux18~6_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux18~1_combout ),
	.datad(\Mux18~8_combout ),
	.cin(gnd),
	.combout(\Mux18~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~9 .lut_mask = 16'hEA62;
defparam \Mux18~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N11
dffeas \my_reg[15][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][13] .is_wysiwyg = "true";
defparam \my_reg[15][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N12
cycloneive_lcell_comb \Mux50~7 (
// Equation(s):
// \Mux50~7_combout  = (dcifimemload_16 & (((\my_reg[13][13]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[12][13]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[12][13]~q ),
	.datab(\my_reg[13][13]~q ),
	.datac(dcifimemload_16),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux50~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~7 .lut_mask = 16'hF0CA;
defparam \Mux50~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N10
cycloneive_lcell_comb \Mux50~8 (
// Equation(s):
// \Mux50~8_combout  = (dcifimemload_17 & ((\Mux50~7_combout  & ((\my_reg[15][13]~q ))) # (!\Mux50~7_combout  & (\my_reg[14][13]~q )))) # (!dcifimemload_17 & (((\Mux50~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[14][13]~q ),
	.datac(\my_reg[15][13]~q ),
	.datad(\Mux50~7_combout ),
	.cin(gnd),
	.combout(\Mux50~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~8 .lut_mask = 16'hF588;
defparam \Mux50~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N7
dffeas \my_reg[3][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][13] .is_wysiwyg = "true";
defparam \my_reg[3][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N6
cycloneive_lcell_comb \Mux50~4 (
// Equation(s):
// \Mux50~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][13]~q ))) # (!dcifimemload_17 & (\my_reg[1][13]~q ))))

	.dataa(\my_reg[1][13]~q ),
	.datab(dcifimemload_17),
	.datac(\my_reg[3][13]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux50~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~4 .lut_mask = 16'hE200;
defparam \Mux50~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N16
cycloneive_lcell_comb \Mux50~5 (
// Equation(s):
// \Mux50~5_combout  = (\Mux50~4_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \my_reg[2][13]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\my_reg[2][13]~q ),
	.datad(\Mux50~4_combout ),
	.cin(gnd),
	.combout(\Mux50~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~5 .lut_mask = 16'hFF40;
defparam \Mux50~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N3
dffeas \my_reg[11][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][13] .is_wysiwyg = "true";
defparam \my_reg[11][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N6
cycloneive_lcell_comb \my_reg[10][13]~feeder (
// Equation(s):
// \my_reg[10][13]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat20),
	.cin(gnd),
	.combout(\my_reg[10][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[10][13]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[10][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y39_N7
dffeas \my_reg[10][13] (
	.clk(CLK),
	.d(\my_reg[10][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][13] .is_wysiwyg = "true";
defparam \my_reg[10][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N24
cycloneive_lcell_comb \Mux50~2 (
// Equation(s):
// \Mux50~2_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\my_reg[10][13]~q )) # (!dcifimemload_17 & ((\my_reg[8][13]~q )))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[10][13]~q ),
	.datac(\my_reg[8][13]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux50~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~2 .lut_mask = 16'hEE50;
defparam \Mux50~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N2
cycloneive_lcell_comb \Mux50~3 (
// Equation(s):
// \Mux50~3_combout  = (dcifimemload_16 & ((\Mux50~2_combout  & ((\my_reg[11][13]~q ))) # (!\Mux50~2_combout  & (\my_reg[9][13]~q )))) # (!dcifimemload_16 & (((\Mux50~2_combout ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[9][13]~q ),
	.datac(\my_reg[11][13]~q ),
	.datad(\Mux50~2_combout ),
	.cin(gnd),
	.combout(\Mux50~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~3 .lut_mask = 16'hF588;
defparam \Mux50~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N16
cycloneive_lcell_comb \Mux50~6 (
// Equation(s):
// \Mux50~6_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\Mux50~3_combout )))) # (!dcifimemload_19 & (!dcifimemload_18 & (\Mux50~5_combout )))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux50~5_combout ),
	.datad(\Mux50~3_combout ),
	.cin(gnd),
	.combout(\Mux50~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~6 .lut_mask = 16'hBA98;
defparam \Mux50~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y32_N11
dffeas \my_reg[5][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][13] .is_wysiwyg = "true";
defparam \my_reg[5][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N10
cycloneive_lcell_comb \Mux50~0 (
// Equation(s):
// \Mux50~0_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][13]~q ))) # (!dcifimemload_16 & (\my_reg[4][13]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[4][13]~q ),
	.datac(\my_reg[5][13]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux50~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~0 .lut_mask = 16'hFA44;
defparam \Mux50~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N4
cycloneive_lcell_comb \Mux50~1 (
// Equation(s):
// \Mux50~1_combout  = (dcifimemload_17 & ((\Mux50~0_combout  & (\my_reg[7][13]~q )) # (!\Mux50~0_combout  & ((\my_reg[6][13]~q ))))) # (!dcifimemload_17 & (((\Mux50~0_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[7][13]~q ),
	.datac(\my_reg[6][13]~q ),
	.datad(\Mux50~0_combout ),
	.cin(gnd),
	.combout(\Mux50~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~1 .lut_mask = 16'hDDA0;
defparam \Mux50~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N14
cycloneive_lcell_comb \my_reg[21][13]~feeder (
// Equation(s):
// \my_reg[21][13]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat20),
	.cin(gnd),
	.combout(\my_reg[21][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][13]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[21][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N15
dffeas \my_reg[21][13] (
	.clk(CLK),
	.d(\my_reg[21][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][13] .is_wysiwyg = "true";
defparam \my_reg[21][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N15
dffeas \my_reg[25][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][13] .is_wysiwyg = "true";
defparam \my_reg[25][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N14
cycloneive_lcell_comb \Mux50~10 (
// Equation(s):
// \Mux50~10_combout  = (dcifimemload_19 & (((\my_reg[25][13]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[17][13]~q  & ((!dcifimemload_18))))

	.dataa(\my_reg[17][13]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[25][13]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux50~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~10 .lut_mask = 16'hCCE2;
defparam \Mux50~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N6
cycloneive_lcell_comb \Mux50~11 (
// Equation(s):
// \Mux50~11_combout  = (dcifimemload_18 & ((\Mux50~10_combout  & ((\my_reg[29][13]~q ))) # (!\Mux50~10_combout  & (\my_reg[21][13]~q )))) # (!dcifimemload_18 & (((\Mux50~10_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[21][13]~q ),
	.datac(\my_reg[29][13]~q ),
	.datad(\Mux50~10_combout ),
	.cin(gnd),
	.combout(\Mux50~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~11 .lut_mask = 16'hF588;
defparam \Mux50~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N26
cycloneive_lcell_comb \my_reg[23][13]~feeder (
// Equation(s):
// \my_reg[23][13]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat20),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[23][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[23][13]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[23][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N27
dffeas \my_reg[23][13] (
	.clk(CLK),
	.d(\my_reg[23][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][13] .is_wysiwyg = "true";
defparam \my_reg[23][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N0
cycloneive_lcell_comb \Mux50~17 (
// Equation(s):
// \Mux50~17_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[27][13]~q ))) # (!dcifimemload_19 & (\my_reg[19][13]~q ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[19][13]~q ),
	.datac(\my_reg[27][13]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux50~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~17 .lut_mask = 16'hFA44;
defparam \Mux50~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N6
cycloneive_lcell_comb \Mux50~18 (
// Equation(s):
// \Mux50~18_combout  = (\Mux50~17_combout  & (((\my_reg[31][13]~q ) # (!dcifimemload_18)))) # (!\Mux50~17_combout  & (\my_reg[23][13]~q  & ((dcifimemload_18))))

	.dataa(\my_reg[23][13]~q ),
	.datab(\my_reg[31][13]~q ),
	.datac(\Mux50~17_combout ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux50~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~18 .lut_mask = 16'hCAF0;
defparam \Mux50~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N8
cycloneive_lcell_comb \my_reg[28][13]~feeder (
// Equation(s):
// \my_reg[28][13]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat20),
	.cin(gnd),
	.combout(\my_reg[28][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[28][13]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[28][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N9
dffeas \my_reg[28][13] (
	.clk(CLK),
	.d(\my_reg[28][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][13] .is_wysiwyg = "true";
defparam \my_reg[28][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N27
dffeas \my_reg[24][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][13] .is_wysiwyg = "true";
defparam \my_reg[24][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N24
cycloneive_lcell_comb \Mux50~14 (
// Equation(s):
// \Mux50~14_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[20][13]~q ))) # (!dcifimemload_18 & (\my_reg[16][13]~q ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[16][13]~q ),
	.datac(\my_reg[20][13]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux50~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~14 .lut_mask = 16'hFA44;
defparam \Mux50~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N26
cycloneive_lcell_comb \Mux50~15 (
// Equation(s):
// \Mux50~15_combout  = (dcifimemload_19 & ((\Mux50~14_combout  & (\my_reg[28][13]~q )) # (!\Mux50~14_combout  & ((\my_reg[24][13]~q ))))) # (!dcifimemload_19 & (((\Mux50~14_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[28][13]~q ),
	.datac(\my_reg[24][13]~q ),
	.datad(\Mux50~14_combout ),
	.cin(gnd),
	.combout(\Mux50~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~15 .lut_mask = 16'hDDA0;
defparam \Mux50~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y42_N9
dffeas \my_reg[22][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][13] .is_wysiwyg = "true";
defparam \my_reg[22][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N8
cycloneive_lcell_comb \Mux50~12 (
// Equation(s):
// \Mux50~12_combout  = (dcifimemload_18 & (((\my_reg[22][13]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[18][13]~q  & ((!dcifimemload_19))))

	.dataa(\my_reg[18][13]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[22][13]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux50~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~12 .lut_mask = 16'hCCE2;
defparam \Mux50~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y42_N31
dffeas \my_reg[26][13] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][13] .is_wysiwyg = "true";
defparam \my_reg[26][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N30
cycloneive_lcell_comb \Mux50~13 (
// Equation(s):
// \Mux50~13_combout  = (\Mux50~12_combout  & ((\my_reg[30][13]~q ) # ((!dcifimemload_19)))) # (!\Mux50~12_combout  & (((\my_reg[26][13]~q  & dcifimemload_19))))

	.dataa(\my_reg[30][13]~q ),
	.datab(\Mux50~12_combout ),
	.datac(\my_reg[26][13]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux50~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~13 .lut_mask = 16'hB8CC;
defparam \Mux50~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N0
cycloneive_lcell_comb \Mux50~16 (
// Equation(s):
// \Mux50~16_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux50~13_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & (\Mux50~15_combout )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux50~15_combout ),
	.datad(\Mux50~13_combout ),
	.cin(gnd),
	.combout(\Mux50~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~16 .lut_mask = 16'hBA98;
defparam \Mux50~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N3
dffeas \my_reg[24][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][12] .is_wysiwyg = "true";
defparam \my_reg[24][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N31
dffeas \my_reg[28][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][12] .is_wysiwyg = "true";
defparam \my_reg[28][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N21
dffeas \my_reg[20][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][12] .is_wysiwyg = "true";
defparam \my_reg[20][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N21
dffeas \my_reg[16][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][12] .is_wysiwyg = "true";
defparam \my_reg[16][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N20
cycloneive_lcell_comb \Mux19~4 (
// Equation(s):
// \Mux19~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[20][12]~q )) # (!dcifimemload_23 & ((\my_reg[16][12]~q )))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[20][12]~q ),
	.datac(\my_reg[16][12]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~4 .lut_mask = 16'hEE50;
defparam \Mux19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N30
cycloneive_lcell_comb \Mux19~5 (
// Equation(s):
// \Mux19~5_combout  = (dcifimemload_24 & ((\Mux19~4_combout  & ((\my_reg[28][12]~q ))) # (!\Mux19~4_combout  & (\my_reg[24][12]~q )))) # (!dcifimemload_24 & (((\Mux19~4_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[24][12]~q ),
	.datac(\my_reg[28][12]~q ),
	.datad(\Mux19~4_combout ),
	.cin(gnd),
	.combout(\Mux19~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~5 .lut_mask = 16'hF588;
defparam \Mux19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N16
cycloneive_lcell_comb \my_reg[30][12]~feeder (
// Equation(s):
// \my_reg[30][12]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat21),
	.cin(gnd),
	.combout(\my_reg[30][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[30][12]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[30][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y29_N17
dffeas \my_reg[30][12] (
	.clk(CLK),
	.d(\my_reg[30][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][12] .is_wysiwyg = "true";
defparam \my_reg[30][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N8
cycloneive_lcell_comb \my_reg[18][12]~feeder (
// Equation(s):
// \my_reg[18][12]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat21),
	.cin(gnd),
	.combout(\my_reg[18][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[18][12]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[18][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y29_N9
dffeas \my_reg[18][12] (
	.clk(CLK),
	.d(\my_reg[18][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][12] .is_wysiwyg = "true";
defparam \my_reg[18][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N18
cycloneive_lcell_comb \Mux19~2 (
// Equation(s):
// \Mux19~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[22][12]~q )) # (!dcifimemload_23 & ((\my_reg[18][12]~q )))))

	.dataa(\my_reg[22][12]~q ),
	.datab(\my_reg[18][12]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~2 .lut_mask = 16'hFA0C;
defparam \Mux19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N6
cycloneive_lcell_comb \Mux19~3 (
// Equation(s):
// \Mux19~3_combout  = (dcifimemload_24 & ((\Mux19~2_combout  & ((\my_reg[30][12]~q ))) # (!\Mux19~2_combout  & (\my_reg[26][12]~q )))) # (!dcifimemload_24 & (((\Mux19~2_combout ))))

	.dataa(\my_reg[26][12]~q ),
	.datab(\my_reg[30][12]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux19~2_combout ),
	.cin(gnd),
	.combout(\Mux19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~3 .lut_mask = 16'hCFA0;
defparam \Mux19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N28
cycloneive_lcell_comb \Mux19~6 (
// Equation(s):
// \Mux19~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux19~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & (\Mux19~5_combout )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux19~5_combout ),
	.datad(\Mux19~3_combout ),
	.cin(gnd),
	.combout(\Mux19~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~6 .lut_mask = 16'hBA98;
defparam \Mux19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N15
dffeas \my_reg[21][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][12] .is_wysiwyg = "true";
defparam \my_reg[21][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N0
cycloneive_lcell_comb \my_reg[25][12]~feeder (
// Equation(s):
// \my_reg[25][12]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat21),
	.cin(gnd),
	.combout(\my_reg[25][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][12]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[25][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y42_N1
dffeas \my_reg[25][12] (
	.clk(CLK),
	.d(\my_reg[25][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][12] .is_wysiwyg = "true";
defparam \my_reg[25][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N20
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\my_reg[25][12]~q ))) # (!dcifimemload_24 & (\my_reg[17][12]~q ))))

	.dataa(\my_reg[17][12]~q ),
	.datab(\my_reg[25][12]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'hFC0A;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N16
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// \Mux19~1_combout  = (\Mux19~0_combout  & ((\my_reg[29][12]~q ) # ((!dcifimemload_23)))) # (!\Mux19~0_combout  & (((\my_reg[21][12]~q  & dcifimemload_23))))

	.dataa(\my_reg[29][12]~q ),
	.datab(\my_reg[21][12]~q ),
	.datac(\Mux19~0_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hACF0;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N2
cycloneive_lcell_comb \my_reg[31][12]~feeder (
// Equation(s):
// \my_reg[31][12]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat21),
	.cin(gnd),
	.combout(\my_reg[31][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[31][12]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[31][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N3
dffeas \my_reg[31][12] (
	.clk(CLK),
	.d(\my_reg[31][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][12] .is_wysiwyg = "true";
defparam \my_reg[31][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N3
dffeas \my_reg[27][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][12] .is_wysiwyg = "true";
defparam \my_reg[27][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N2
cycloneive_lcell_comb \Mux19~7 (
// Equation(s):
// \Mux19~7_combout  = (dcifimemload_24 & (((\my_reg[27][12]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\my_reg[19][12]~q  & ((!dcifimemload_23))))

	.dataa(\my_reg[19][12]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[27][12]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux19~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~7 .lut_mask = 16'hCCE2;
defparam \Mux19~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N12
cycloneive_lcell_comb \Mux19~8 (
// Equation(s):
// \Mux19~8_combout  = (dcifimemload_23 & ((\Mux19~7_combout  & ((\my_reg[31][12]~q ))) # (!\Mux19~7_combout  & (\my_reg[23][12]~q )))) # (!dcifimemload_23 & (((\Mux19~7_combout ))))

	.dataa(\my_reg[23][12]~q ),
	.datab(\my_reg[31][12]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux19~7_combout ),
	.cin(gnd),
	.combout(\Mux19~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~8 .lut_mask = 16'hCFA0;
defparam \Mux19~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N22
cycloneive_lcell_comb \Mux19~9 (
// Equation(s):
// \Mux19~9_combout  = (dcifimemload_21 & ((\Mux19~6_combout  & ((\Mux19~8_combout ))) # (!\Mux19~6_combout  & (\Mux19~1_combout )))) # (!dcifimemload_21 & (\Mux19~6_combout ))

	.dataa(dcifimemload_21),
	.datab(\Mux19~6_combout ),
	.datac(\Mux19~1_combout ),
	.datad(\Mux19~8_combout ),
	.cin(gnd),
	.combout(\Mux19~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~9 .lut_mask = 16'hEC64;
defparam \Mux19~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N25
dffeas \my_reg[1][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][12] .is_wysiwyg = "true";
defparam \my_reg[1][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N10
cycloneive_lcell_comb \Mux19~14 (
// Equation(s):
// \Mux19~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & (\my_reg[3][12]~q )) # (!dcifimemload_22 & ((\my_reg[1][12]~q )))))

	.dataa(\my_reg[3][12]~q ),
	.datab(dcifimemload_21),
	.datac(dcifimemload_22),
	.datad(\my_reg[1][12]~q ),
	.cin(gnd),
	.combout(\Mux19~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~14 .lut_mask = 16'h8C80;
defparam \Mux19~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N26
cycloneive_lcell_comb \Mux19~15 (
// Equation(s):
// \Mux19~15_combout  = (\Mux19~14_combout ) # ((\my_reg[2][12]~q  & (!dcifimemload_21 & dcifimemload_22)))

	.dataa(\my_reg[2][12]~q ),
	.datab(dcifimemload_21),
	.datac(dcifimemload_22),
	.datad(\Mux19~14_combout ),
	.cin(gnd),
	.combout(\Mux19~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~15 .lut_mask = 16'hFF20;
defparam \Mux19~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y30_N5
dffeas \my_reg[9][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][12] .is_wysiwyg = "true";
defparam \my_reg[9][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N27
dffeas \my_reg[11][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][12] .is_wysiwyg = "true";
defparam \my_reg[11][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N2
cycloneive_lcell_comb \my_reg[8][12]~feeder (
// Equation(s):
// \my_reg[8][12]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat21),
	.cin(gnd),
	.combout(\my_reg[8][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[8][12]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[8][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N3
dffeas \my_reg[8][12] (
	.clk(CLK),
	.d(\my_reg[8][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][12] .is_wysiwyg = "true";
defparam \my_reg[8][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N28
cycloneive_lcell_comb \Mux19~12 (
// Equation(s):
// \Mux19~12_combout  = (dcifimemload_22 & ((\my_reg[10][12]~q ) # ((dcifimemload_21)))) # (!dcifimemload_22 & (((\my_reg[8][12]~q  & !dcifimemload_21))))

	.dataa(\my_reg[10][12]~q ),
	.datab(\my_reg[8][12]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux19~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~12 .lut_mask = 16'hF0AC;
defparam \Mux19~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N26
cycloneive_lcell_comb \Mux19~13 (
// Equation(s):
// \Mux19~13_combout  = (dcifimemload_21 & ((\Mux19~12_combout  & ((\my_reg[11][12]~q ))) # (!\Mux19~12_combout  & (\my_reg[9][12]~q )))) # (!dcifimemload_21 & (((\Mux19~12_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][12]~q ),
	.datac(\my_reg[11][12]~q ),
	.datad(\Mux19~12_combout ),
	.cin(gnd),
	.combout(\Mux19~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~13 .lut_mask = 16'hF588;
defparam \Mux19~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N16
cycloneive_lcell_comb \Mux19~16 (
// Equation(s):
// \Mux19~16_combout  = (dcifimemload_23 & (dcifimemload_24)) # (!dcifimemload_23 & ((dcifimemload_24 & ((\Mux19~13_combout ))) # (!dcifimemload_24 & (\Mux19~15_combout ))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux19~15_combout ),
	.datad(\Mux19~13_combout ),
	.cin(gnd),
	.combout(\Mux19~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~16 .lut_mask = 16'hDC98;
defparam \Mux19~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N8
cycloneive_lcell_comb \my_reg[12][12]~feeder (
// Equation(s):
// \my_reg[12][12]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat21),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[12][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[12][12]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[12][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N9
dffeas \my_reg[12][12] (
	.clk(CLK),
	.d(\my_reg[12][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][12] .is_wysiwyg = "true";
defparam \my_reg[12][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N27
dffeas \my_reg[13][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][12] .is_wysiwyg = "true";
defparam \my_reg[13][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N26
cycloneive_lcell_comb \Mux19~17 (
// Equation(s):
// \Mux19~17_combout  = (dcifimemload_21 & (((\my_reg[13][12]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\my_reg[12][12]~q  & ((!dcifimemload_22))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[12][12]~q ),
	.datac(\my_reg[13][12]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux19~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~17 .lut_mask = 16'hAAE4;
defparam \Mux19~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N13
dffeas \my_reg[14][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][12] .is_wysiwyg = "true";
defparam \my_reg[14][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N30
cycloneive_lcell_comb \Mux19~18 (
// Equation(s):
// \Mux19~18_combout  = (dcifimemload_22 & ((\Mux19~17_combout  & (\my_reg[15][12]~q )) # (!\Mux19~17_combout  & ((\my_reg[14][12]~q ))))) # (!dcifimemload_22 & (((\Mux19~17_combout ))))

	.dataa(\my_reg[15][12]~q ),
	.datab(dcifimemload_22),
	.datac(\Mux19~17_combout ),
	.datad(\my_reg[14][12]~q ),
	.cin(gnd),
	.combout(\Mux19~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~18 .lut_mask = 16'hBCB0;
defparam \Mux19~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N28
cycloneive_lcell_comb \my_reg[6][12]~feeder (
// Equation(s):
// \my_reg[6][12]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat21),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[6][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[6][12]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[6][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y43_N29
dffeas \my_reg[6][12] (
	.clk(CLK),
	.d(\my_reg[6][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][12] .is_wysiwyg = "true";
defparam \my_reg[6][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N29
dffeas \my_reg[4][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][12] .is_wysiwyg = "true";
defparam \my_reg[4][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N8
cycloneive_lcell_comb \Mux19~10 (
// Equation(s):
// \Mux19~10_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\my_reg[5][12]~q )) # (!dcifimemload_21 & ((\my_reg[4][12]~q )))))

	.dataa(\my_reg[5][12]~q ),
	.datab(\my_reg[4][12]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux19~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~10 .lut_mask = 16'hFA0C;
defparam \Mux19~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N15
dffeas \my_reg[7][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][12] .is_wysiwyg = "true";
defparam \my_reg[7][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N26
cycloneive_lcell_comb \Mux19~11 (
// Equation(s):
// \Mux19~11_combout  = (dcifimemload_22 & ((\Mux19~10_combout  & ((\my_reg[7][12]~q ))) # (!\Mux19~10_combout  & (\my_reg[6][12]~q )))) # (!dcifimemload_22 & (((\Mux19~10_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[6][12]~q ),
	.datac(\Mux19~10_combout ),
	.datad(\my_reg[7][12]~q ),
	.cin(gnd),
	.combout(\Mux19~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~11 .lut_mask = 16'hF858;
defparam \Mux19~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N0
cycloneive_lcell_comb \Mux19~19 (
// Equation(s):
// \Mux19~19_combout  = (dcifimemload_23 & ((\Mux19~16_combout  & (\Mux19~18_combout )) # (!\Mux19~16_combout  & ((\Mux19~11_combout ))))) # (!dcifimemload_23 & (\Mux19~16_combout ))

	.dataa(dcifimemload_23),
	.datab(\Mux19~16_combout ),
	.datac(\Mux19~18_combout ),
	.datad(\Mux19~11_combout ),
	.cin(gnd),
	.combout(\Mux19~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~19 .lut_mask = 16'hE6C4;
defparam \Mux19~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y30_N11
dffeas \my_reg[10][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][12] .is_wysiwyg = "true";
defparam \my_reg[10][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N10
cycloneive_lcell_comb \Mux51~0 (
// Equation(s):
// \Mux51~0_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[10][12]~q ))) # (!dcifimemload_17 & (\my_reg[8][12]~q ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[8][12]~q ),
	.datac(\my_reg[10][12]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux51~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~0 .lut_mask = 16'hFA44;
defparam \Mux51~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N4
cycloneive_lcell_comb \Mux51~1 (
// Equation(s):
// \Mux51~1_combout  = (dcifimemload_16 & ((\Mux51~0_combout  & (\my_reg[11][12]~q )) # (!\Mux51~0_combout  & ((\my_reg[9][12]~q ))))) # (!dcifimemload_16 & (((\Mux51~0_combout ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[11][12]~q ),
	.datac(\my_reg[9][12]~q ),
	.datad(\Mux51~0_combout ),
	.cin(gnd),
	.combout(\Mux51~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~1 .lut_mask = 16'hDDA0;
defparam \Mux51~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N23
dffeas \my_reg[15][12] (
	.clk(CLK),
	.d(wdat21),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][12] .is_wysiwyg = "true";
defparam \my_reg[15][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N30
cycloneive_lcell_comb \Mux51~7 (
// Equation(s):
// \Mux51~7_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\my_reg[13][12]~q )) # (!dcifimemload_16 & ((\my_reg[12][12]~q )))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[13][12]~q ),
	.datac(\my_reg[12][12]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux51~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~7 .lut_mask = 16'hEE50;
defparam \Mux51~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N12
cycloneive_lcell_comb \Mux51~8 (
// Equation(s):
// \Mux51~8_combout  = (\Mux51~7_combout  & ((\my_reg[15][12]~q ) # ((!dcifimemload_17)))) # (!\Mux51~7_combout  & (((\my_reg[14][12]~q  & dcifimemload_17))))

	.dataa(\my_reg[15][12]~q ),
	.datab(\Mux51~7_combout ),
	.datac(\my_reg[14][12]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux51~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~8 .lut_mask = 16'hB8CC;
defparam \Mux51~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N28
cycloneive_lcell_comb \Mux51~2 (
// Equation(s):
// \Mux51~2_combout  = (dcifimemload_16 & ((\my_reg[5][12]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\my_reg[4][12]~q  & !dcifimemload_17))))

	.dataa(\my_reg[5][12]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[4][12]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux51~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~2 .lut_mask = 16'hCCB8;
defparam \Mux51~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N14
cycloneive_lcell_comb \Mux51~3 (
// Equation(s):
// \Mux51~3_combout  = (dcifimemload_17 & ((\Mux51~2_combout  & ((\my_reg[7][12]~q ))) # (!\Mux51~2_combout  & (\my_reg[6][12]~q )))) # (!dcifimemload_17 & (((\Mux51~2_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[6][12]~q ),
	.datac(\my_reg[7][12]~q ),
	.datad(\Mux51~2_combout ),
	.cin(gnd),
	.combout(\Mux51~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~3 .lut_mask = 16'hF588;
defparam \Mux51~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N13
dffeas \my_reg[2][12] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][12] .is_wysiwyg = "true";
defparam \my_reg[2][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N26
cycloneive_lcell_comb \my_reg[3][12]~feeder (
// Equation(s):
// \my_reg[3][12]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat21),
	.cin(gnd),
	.combout(\my_reg[3][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[3][12]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[3][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y37_N27
dffeas \my_reg[3][12] (
	.clk(CLK),
	.d(\my_reg[3][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][12] .is_wysiwyg = "true";
defparam \my_reg[3][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N24
cycloneive_lcell_comb \Mux51~4 (
// Equation(s):
// \Mux51~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\my_reg[3][12]~q )) # (!dcifimemload_17 & ((\my_reg[1][12]~q )))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[3][12]~q ),
	.datac(\my_reg[1][12]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux51~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~4 .lut_mask = 16'hD800;
defparam \Mux51~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N12
cycloneive_lcell_comb \Mux51~5 (
// Equation(s):
// \Mux51~5_combout  = (\Mux51~4_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \my_reg[2][12]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\my_reg[2][12]~q ),
	.datad(\Mux51~4_combout ),
	.cin(gnd),
	.combout(\Mux51~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~5 .lut_mask = 16'hFF20;
defparam \Mux51~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N20
cycloneive_lcell_comb \Mux51~6 (
// Equation(s):
// \Mux51~6_combout  = (dcifimemload_18 & ((dcifimemload_19) # ((\Mux51~3_combout )))) # (!dcifimemload_18 & (!dcifimemload_19 & ((\Mux51~5_combout ))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux51~3_combout ),
	.datad(\Mux51~5_combout ),
	.cin(gnd),
	.combout(\Mux51~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~6 .lut_mask = 16'hB9A8;
defparam \Mux51~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N14
cycloneive_lcell_comb \Mux51~10 (
// Equation(s):
// \Mux51~10_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[21][12]~q ))) # (!dcifimemload_18 & (\my_reg[17][12]~q ))))

	.dataa(\my_reg[17][12]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[21][12]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux51~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~10 .lut_mask = 16'hFC22;
defparam \Mux51~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N22
cycloneive_lcell_comb \my_reg[29][12]~feeder (
// Equation(s):
// \my_reg[29][12]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat21),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[29][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[29][12]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[29][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N23
dffeas \my_reg[29][12] (
	.clk(CLK),
	.d(\my_reg[29][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][12] .is_wysiwyg = "true";
defparam \my_reg[29][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N2
cycloneive_lcell_comb \Mux51~11 (
// Equation(s):
// \Mux51~11_combout  = (\Mux51~10_combout  & (((\my_reg[29][12]~q ) # (!dcifimemload_19)))) # (!\Mux51~10_combout  & (\my_reg[25][12]~q  & ((dcifimemload_19))))

	.dataa(\Mux51~10_combout ),
	.datab(\my_reg[25][12]~q ),
	.datac(\my_reg[29][12]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux51~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~11 .lut_mask = 16'hE4AA;
defparam \Mux51~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N16
cycloneive_lcell_comb \my_reg[19][12]~feeder (
// Equation(s):
// \my_reg[19][12]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat21),
	.cin(gnd),
	.combout(\my_reg[19][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[19][12]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[19][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y34_N17
dffeas \my_reg[19][12] (
	.clk(CLK),
	.d(\my_reg[19][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][12] .is_wysiwyg = "true";
defparam \my_reg[19][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N10
cycloneive_lcell_comb \Mux51~17 (
// Equation(s):
// \Mux51~17_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\my_reg[23][12]~q )) # (!dcifimemload_18 & ((\my_reg[19][12]~q )))))

	.dataa(\my_reg[23][12]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[19][12]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux51~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~17 .lut_mask = 16'hEE30;
defparam \Mux51~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N24
cycloneive_lcell_comb \Mux51~18 (
// Equation(s):
// \Mux51~18_combout  = (dcifimemload_19 & ((\Mux51~17_combout  & ((\my_reg[31][12]~q ))) # (!\Mux51~17_combout  & (\my_reg[27][12]~q )))) # (!dcifimemload_19 & (((\Mux51~17_combout ))))

	.dataa(\my_reg[27][12]~q ),
	.datab(\my_reg[31][12]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux51~17_combout ),
	.cin(gnd),
	.combout(\Mux51~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~18 .lut_mask = 16'hCFA0;
defparam \Mux51~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N2
cycloneive_lcell_comb \Mux51~14 (
// Equation(s):
// \Mux51~14_combout  = (dcifimemload_19 & (((\my_reg[24][12]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[16][12]~q  & ((!dcifimemload_18))))

	.dataa(\my_reg[16][12]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[24][12]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux51~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~14 .lut_mask = 16'hCCE2;
defparam \Mux51~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N20
cycloneive_lcell_comb \Mux51~15 (
// Equation(s):
// \Mux51~15_combout  = (dcifimemload_18 & ((\Mux51~14_combout  & (\my_reg[28][12]~q )) # (!\Mux51~14_combout  & ((\my_reg[20][12]~q ))))) # (!dcifimemload_18 & (((\Mux51~14_combout ))))

	.dataa(\my_reg[28][12]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[20][12]~q ),
	.datad(\Mux51~14_combout ),
	.cin(gnd),
	.combout(\Mux51~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~15 .lut_mask = 16'hBBC0;
defparam \Mux51~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N4
cycloneive_lcell_comb \my_reg[26][12]~feeder (
// Equation(s):
// \my_reg[26][12]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat21),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[26][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[26][12]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[26][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y29_N5
dffeas \my_reg[26][12] (
	.clk(CLK),
	.d(\my_reg[26][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][12] .is_wysiwyg = "true";
defparam \my_reg[26][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N28
cycloneive_lcell_comb \Mux51~12 (
// Equation(s):
// \Mux51~12_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[26][12]~q ))) # (!dcifimemload_19 & (\my_reg[18][12]~q ))))

	.dataa(\my_reg[18][12]~q ),
	.datab(\my_reg[26][12]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux51~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~12 .lut_mask = 16'hFC0A;
defparam \Mux51~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N14
cycloneive_lcell_comb \Mux51~13 (
// Equation(s):
// \Mux51~13_combout  = (dcifimemload_18 & ((\Mux51~12_combout  & ((\my_reg[30][12]~q ))) # (!\Mux51~12_combout  & (\my_reg[22][12]~q )))) # (!dcifimemload_18 & (((\Mux51~12_combout ))))

	.dataa(\my_reg[22][12]~q ),
	.datab(\my_reg[30][12]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux51~12_combout ),
	.cin(gnd),
	.combout(\Mux51~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~13 .lut_mask = 16'hCFA0;
defparam \Mux51~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N14
cycloneive_lcell_comb \Mux51~16 (
// Equation(s):
// \Mux51~16_combout  = (dcifimemload_17 & (((dcifimemload_16) # (\Mux51~13_combout )))) # (!dcifimemload_17 & (\Mux51~15_combout  & (!dcifimemload_16)))

	.dataa(dcifimemload_17),
	.datab(\Mux51~15_combout ),
	.datac(dcifimemload_16),
	.datad(\Mux51~13_combout ),
	.cin(gnd),
	.combout(\Mux51~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~16 .lut_mask = 16'hAEA4;
defparam \Mux51~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N15
dffeas \my_reg[7][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][11] .is_wysiwyg = "true";
defparam \my_reg[7][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N29
dffeas \my_reg[4][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][11] .is_wysiwyg = "true";
defparam \my_reg[4][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N28
cycloneive_lcell_comb \Mux20~12 (
// Equation(s):
// \Mux20~12_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\my_reg[5][11]~q )) # (!dcifimemload_21 & ((\my_reg[4][11]~q )))))

	.dataa(\my_reg[5][11]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[4][11]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux20~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~12 .lut_mask = 16'hEE30;
defparam \Mux20~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N14
cycloneive_lcell_comb \Mux20~13 (
// Equation(s):
// \Mux20~13_combout  = (dcifimemload_22 & ((\Mux20~12_combout  & ((\my_reg[7][11]~q ))) # (!\Mux20~12_combout  & (\my_reg[6][11]~q )))) # (!dcifimemload_22 & (((\Mux20~12_combout ))))

	.dataa(\my_reg[6][11]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[7][11]~q ),
	.datad(\Mux20~12_combout ),
	.cin(gnd),
	.combout(\Mux20~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~13 .lut_mask = 16'hF388;
defparam \Mux20~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N7
dffeas \my_reg[1][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][11] .is_wysiwyg = "true";
defparam \my_reg[1][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N21
dffeas \my_reg[3][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][11] .is_wysiwyg = "true";
defparam \my_reg[3][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N20
cycloneive_lcell_comb \Mux20~14 (
// Equation(s):
// \Mux20~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][11]~q ))) # (!dcifimemload_22 & (\my_reg[1][11]~q ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[1][11]~q ),
	.datac(\my_reg[3][11]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux20~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~14 .lut_mask = 16'hA088;
defparam \Mux20~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N10
cycloneive_lcell_comb \Mux20~15 (
// Equation(s):
// \Mux20~15_combout  = (\Mux20~14_combout ) # ((\my_reg[2][11]~q  & (dcifimemload_22 & !dcifimemload_21)))

	.dataa(\my_reg[2][11]~q ),
	.datab(dcifimemload_22),
	.datac(dcifimemload_21),
	.datad(\Mux20~14_combout ),
	.cin(gnd),
	.combout(\Mux20~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~15 .lut_mask = 16'hFF08;
defparam \Mux20~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N16
cycloneive_lcell_comb \Mux20~16 (
// Equation(s):
// \Mux20~16_combout  = (dcifimemload_23 & ((dcifimemload_24) # ((\Mux20~13_combout )))) # (!dcifimemload_23 & (!dcifimemload_24 & ((\Mux20~15_combout ))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux20~13_combout ),
	.datad(\Mux20~15_combout ),
	.cin(gnd),
	.combout(\Mux20~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~16 .lut_mask = 16'hB9A8;
defparam \Mux20~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N21
dffeas \my_reg[14][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][11] .is_wysiwyg = "true";
defparam \my_reg[14][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N25
dffeas \my_reg[13][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][11] .is_wysiwyg = "true";
defparam \my_reg[13][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N24
cycloneive_lcell_comb \Mux20~17 (
// Equation(s):
// \Mux20~17_combout  = (dcifimemload_21 & (((\my_reg[13][11]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\my_reg[12][11]~q  & ((!dcifimemload_22))))

	.dataa(\my_reg[12][11]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[13][11]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux20~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~17 .lut_mask = 16'hCCE2;
defparam \Mux20~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N22
cycloneive_lcell_comb \Mux20~18 (
// Equation(s):
// \Mux20~18_combout  = (dcifimemload_22 & ((\Mux20~17_combout  & (\my_reg[15][11]~q )) # (!\Mux20~17_combout  & ((\my_reg[14][11]~q ))))) # (!dcifimemload_22 & (((\Mux20~17_combout ))))

	.dataa(\my_reg[15][11]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[14][11]~q ),
	.datad(\Mux20~17_combout ),
	.cin(gnd),
	.combout(\Mux20~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~18 .lut_mask = 16'hBBC0;
defparam \Mux20~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N27
dffeas \my_reg[11][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][11] .is_wysiwyg = "true";
defparam \my_reg[11][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N27
dffeas \my_reg[10][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][11] .is_wysiwyg = "true";
defparam \my_reg[10][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N26
cycloneive_lcell_comb \Mux20~10 (
// Equation(s):
// \Mux20~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[10][11]~q ))) # (!dcifimemload_22 & (\my_reg[8][11]~q ))))

	.dataa(\my_reg[8][11]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[10][11]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux20~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~10 .lut_mask = 16'hFC22;
defparam \Mux20~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N16
cycloneive_lcell_comb \Mux20~11 (
// Equation(s):
// \Mux20~11_combout  = (\Mux20~10_combout  & (((\my_reg[11][11]~q ) # (!dcifimemload_21)))) # (!\Mux20~10_combout  & (\my_reg[9][11]~q  & ((dcifimemload_21))))

	.dataa(\my_reg[9][11]~q ),
	.datab(\my_reg[11][11]~q ),
	.datac(\Mux20~10_combout ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux20~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~11 .lut_mask = 16'hCAF0;
defparam \Mux20~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N8
cycloneive_lcell_comb \Mux20~19 (
// Equation(s):
// \Mux20~19_combout  = (dcifimemload_24 & ((\Mux20~16_combout  & (\Mux20~18_combout )) # (!\Mux20~16_combout  & ((\Mux20~11_combout ))))) # (!dcifimemload_24 & (\Mux20~16_combout ))

	.dataa(dcifimemload_24),
	.datab(\Mux20~16_combout ),
	.datac(\Mux20~18_combout ),
	.datad(\Mux20~11_combout ),
	.cin(gnd),
	.combout(\Mux20~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~19 .lut_mask = 16'hE6C4;
defparam \Mux20~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N27
dffeas \my_reg[31][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][11] .is_wysiwyg = "true";
defparam \my_reg[31][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N19
dffeas \my_reg[19][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][11] .is_wysiwyg = "true";
defparam \my_reg[19][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N18
cycloneive_lcell_comb \Mux20~7 (
// Equation(s):
// \Mux20~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[23][11]~q )) # (!dcifimemload_23 & ((\my_reg[19][11]~q )))))

	.dataa(\my_reg[23][11]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[19][11]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux20~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~7 .lut_mask = 16'hEE30;
defparam \Mux20~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N26
cycloneive_lcell_comb \Mux20~8 (
// Equation(s):
// \Mux20~8_combout  = (dcifimemload_24 & ((\Mux20~7_combout  & ((\my_reg[31][11]~q ))) # (!\Mux20~7_combout  & (\my_reg[27][11]~q )))) # (!dcifimemload_24 & (((\Mux20~7_combout ))))

	.dataa(\my_reg[27][11]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[31][11]~q ),
	.datad(\Mux20~7_combout ),
	.cin(gnd),
	.combout(\Mux20~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~8 .lut_mask = 16'hF388;
defparam \Mux20~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y37_N21
dffeas \my_reg[20][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][11] .is_wysiwyg = "true";
defparam \my_reg[20][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N27
dffeas \my_reg[28][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][11] .is_wysiwyg = "true";
defparam \my_reg[28][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N27
dffeas \my_reg[24][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][11] .is_wysiwyg = "true";
defparam \my_reg[24][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N1
dffeas \my_reg[16][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][11] .is_wysiwyg = "true";
defparam \my_reg[16][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N0
cycloneive_lcell_comb \Mux20~4 (
// Equation(s):
// \Mux20~4_combout  = (dcifimemload_24 & ((\my_reg[24][11]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\my_reg[16][11]~q  & !dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[24][11]~q ),
	.datac(\my_reg[16][11]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~4 .lut_mask = 16'hAAD8;
defparam \Mux20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N26
cycloneive_lcell_comb \Mux20~5 (
// Equation(s):
// \Mux20~5_combout  = (dcifimemload_23 & ((\Mux20~4_combout  & ((\my_reg[28][11]~q ))) # (!\Mux20~4_combout  & (\my_reg[20][11]~q )))) # (!dcifimemload_23 & (((\Mux20~4_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[20][11]~q ),
	.datac(\my_reg[28][11]~q ),
	.datad(\Mux20~4_combout ),
	.cin(gnd),
	.combout(\Mux20~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~5 .lut_mask = 16'hF588;
defparam \Mux20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N17
dffeas \my_reg[30][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][11] .is_wysiwyg = "true";
defparam \my_reg[30][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N30
cycloneive_lcell_comb \my_reg[18][11]~feeder (
// Equation(s):
// \my_reg[18][11]~feeder_combout  = \wdat~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat22),
	.cin(gnd),
	.combout(\my_reg[18][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[18][11]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[18][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N31
dffeas \my_reg[18][11] (
	.clk(CLK),
	.d(\my_reg[18][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][11] .is_wysiwyg = "true";
defparam \my_reg[18][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N20
cycloneive_lcell_comb \Mux20~2 (
// Equation(s):
// \Mux20~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[26][11]~q )) # (!dcifimemload_24 & ((\my_reg[18][11]~q )))))

	.dataa(\my_reg[26][11]~q ),
	.datab(\my_reg[18][11]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux20~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~2 .lut_mask = 16'hFA0C;
defparam \Mux20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N22
cycloneive_lcell_comb \Mux20~3 (
// Equation(s):
// \Mux20~3_combout  = (dcifimemload_23 & ((\Mux20~2_combout  & ((\my_reg[30][11]~q ))) # (!\Mux20~2_combout  & (\my_reg[22][11]~q )))) # (!dcifimemload_23 & (((\Mux20~2_combout ))))

	.dataa(\my_reg[22][11]~q ),
	.datab(\my_reg[30][11]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux20~2_combout ),
	.cin(gnd),
	.combout(\Mux20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~3 .lut_mask = 16'hCFA0;
defparam \Mux20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N26
cycloneive_lcell_comb \Mux20~6 (
// Equation(s):
// \Mux20~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux20~3_combout ))) # (!dcifimemload_22 & (\Mux20~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux20~5_combout ),
	.datad(\Mux20~3_combout ),
	.cin(gnd),
	.combout(\Mux20~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~6 .lut_mask = 16'hDC98;
defparam \Mux20~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N21
dffeas \my_reg[29][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][11] .is_wysiwyg = "true";
defparam \my_reg[29][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N13
dffeas \my_reg[17][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][11] .is_wysiwyg = "true";
defparam \my_reg[17][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N12
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (dcifimemload_23 & ((\my_reg[21][11]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[17][11]~q  & !dcifimemload_24))))

	.dataa(\my_reg[21][11]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[17][11]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'hCCB8;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N20
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// \Mux20~1_combout  = (dcifimemload_24 & ((\Mux20~0_combout  & ((\my_reg[29][11]~q ))) # (!\Mux20~0_combout  & (\my_reg[25][11]~q )))) # (!dcifimemload_24 & (((\Mux20~0_combout ))))

	.dataa(\my_reg[25][11]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[29][11]~q ),
	.datad(\Mux20~0_combout ),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'hF388;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N28
cycloneive_lcell_comb \Mux20~9 (
// Equation(s):
// \Mux20~9_combout  = (dcifimemload_21 & ((\Mux20~6_combout  & (\Mux20~8_combout )) # (!\Mux20~6_combout  & ((\Mux20~1_combout ))))) # (!dcifimemload_21 & (((\Mux20~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux20~8_combout ),
	.datac(\Mux20~6_combout ),
	.datad(\Mux20~1_combout ),
	.cin(gnd),
	.combout(\Mux20~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~9 .lut_mask = 16'hDAD0;
defparam \Mux20~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N3
dffeas \my_reg[12][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][11] .is_wysiwyg = "true";
defparam \my_reg[12][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N2
cycloneive_lcell_comb \Mux52~7 (
// Equation(s):
// \Mux52~7_combout  = (dcifimemload_16 & ((\my_reg[13][11]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\my_reg[12][11]~q  & !dcifimemload_17))))

	.dataa(\my_reg[13][11]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[12][11]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux52~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~7 .lut_mask = 16'hCCB8;
defparam \Mux52~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N5
dffeas \my_reg[15][11] (
	.clk(CLK),
	.d(wdat22),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][11] .is_wysiwyg = "true";
defparam \my_reg[15][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N20
cycloneive_lcell_comb \Mux52~8 (
// Equation(s):
// \Mux52~8_combout  = (dcifimemload_17 & ((\Mux52~7_combout  & ((\my_reg[15][11]~q ))) # (!\Mux52~7_combout  & (\my_reg[14][11]~q )))) # (!dcifimemload_17 & (\Mux52~7_combout ))

	.dataa(dcifimemload_17),
	.datab(\Mux52~7_combout ),
	.datac(\my_reg[14][11]~q ),
	.datad(\my_reg[15][11]~q ),
	.cin(gnd),
	.combout(\Mux52~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~8 .lut_mask = 16'hEC64;
defparam \Mux52~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N26
cycloneive_lcell_comb \my_reg[9][11]~feeder (
// Equation(s):
// \my_reg[9][11]~feeder_combout  = \wdat~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat22),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[9][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[9][11]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[9][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N27
dffeas \my_reg[9][11] (
	.clk(CLK),
	.d(\my_reg[9][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][11] .is_wysiwyg = "true";
defparam \my_reg[9][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N21
dffeas \my_reg[8][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][11] .is_wysiwyg = "true";
defparam \my_reg[8][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N20
cycloneive_lcell_comb \Mux52~2 (
// Equation(s):
// \Mux52~2_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\my_reg[10][11]~q )) # (!dcifimemload_17 & ((\my_reg[8][11]~q )))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[10][11]~q ),
	.datac(\my_reg[8][11]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux52~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~2 .lut_mask = 16'hEE50;
defparam \Mux52~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N26
cycloneive_lcell_comb \Mux52~3 (
// Equation(s):
// \Mux52~3_combout  = (dcifimemload_16 & ((\Mux52~2_combout  & ((\my_reg[11][11]~q ))) # (!\Mux52~2_combout  & (\my_reg[9][11]~q )))) # (!dcifimemload_16 & (((\Mux52~2_combout ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[9][11]~q ),
	.datac(\my_reg[11][11]~q ),
	.datad(\Mux52~2_combout ),
	.cin(gnd),
	.combout(\Mux52~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~3 .lut_mask = 16'hF588;
defparam \Mux52~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N13
dffeas \my_reg[2][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][11] .is_wysiwyg = "true";
defparam \my_reg[2][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N12
cycloneive_lcell_comb \Mux52~5 (
// Equation(s):
// \Mux52~5_combout  = (\Mux52~4_combout ) # ((!dcifimemload_16 & (\my_reg[2][11]~q  & dcifimemload_17)))

	.dataa(\Mux52~4_combout ),
	.datab(dcifimemload_16),
	.datac(\my_reg[2][11]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux52~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~5 .lut_mask = 16'hBAAA;
defparam \Mux52~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N8
cycloneive_lcell_comb \Mux52~6 (
// Equation(s):
// \Mux52~6_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & (\Mux52~3_combout )) # (!dcifimemload_19 & ((\Mux52~5_combout )))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux52~3_combout ),
	.datad(\Mux52~5_combout ),
	.cin(gnd),
	.combout(\Mux52~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~6 .lut_mask = 16'hD9C8;
defparam \Mux52~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y32_N1
dffeas \my_reg[6][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][11] .is_wysiwyg = "true";
defparam \my_reg[6][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y32_N19
dffeas \my_reg[5][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][11] .is_wysiwyg = "true";
defparam \my_reg[5][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N18
cycloneive_lcell_comb \Mux52~0 (
// Equation(s):
// \Mux52~0_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][11]~q ))) # (!dcifimemload_16 & (\my_reg[4][11]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[4][11]~q ),
	.datac(\my_reg[5][11]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux52~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~0 .lut_mask = 16'hFA44;
defparam \Mux52~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N0
cycloneive_lcell_comb \Mux52~1 (
// Equation(s):
// \Mux52~1_combout  = (dcifimemload_17 & ((\Mux52~0_combout  & (\my_reg[7][11]~q )) # (!\Mux52~0_combout  & ((\my_reg[6][11]~q ))))) # (!dcifimemload_17 & (((\Mux52~0_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[7][11]~q ),
	.datac(\my_reg[6][11]~q ),
	.datad(\Mux52~0_combout ),
	.cin(gnd),
	.combout(\Mux52~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~1 .lut_mask = 16'hDDA0;
defparam \Mux52~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N6
cycloneive_lcell_comb \my_reg[27][11]~feeder (
// Equation(s):
// \my_reg[27][11]~feeder_combout  = \wdat~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat22),
	.cin(gnd),
	.combout(\my_reg[27][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[27][11]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[27][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y32_N7
dffeas \my_reg[27][11] (
	.clk(CLK),
	.d(\my_reg[27][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][11] .is_wysiwyg = "true";
defparam \my_reg[27][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N8
cycloneive_lcell_comb \Mux52~17 (
// Equation(s):
// \Mux52~17_combout  = (dcifimemload_19 & (((\my_reg[27][11]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[19][11]~q  & ((!dcifimemload_18))))

	.dataa(\my_reg[19][11]~q ),
	.datab(\my_reg[27][11]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux52~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~17 .lut_mask = 16'hF0CA;
defparam \Mux52~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N1
dffeas \my_reg[23][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][11] .is_wysiwyg = "true";
defparam \my_reg[23][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N0
cycloneive_lcell_comb \Mux52~18 (
// Equation(s):
// \Mux52~18_combout  = (\Mux52~17_combout  & ((\my_reg[31][11]~q ) # ((!dcifimemload_18)))) # (!\Mux52~17_combout  & (((\my_reg[23][11]~q  & dcifimemload_18))))

	.dataa(\my_reg[31][11]~q ),
	.datab(\Mux52~17_combout ),
	.datac(\my_reg[23][11]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux52~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~18 .lut_mask = 16'hB8CC;
defparam \Mux52~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N12
cycloneive_lcell_comb \my_reg[21][11]~feeder (
// Equation(s):
// \my_reg[21][11]~feeder_combout  = \wdat~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat22),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[21][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][11]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[21][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N13
dffeas \my_reg[21][11] (
	.clk(CLK),
	.d(\my_reg[21][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][11] .is_wysiwyg = "true";
defparam \my_reg[21][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N11
dffeas \my_reg[25][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][11] .is_wysiwyg = "true";
defparam \my_reg[25][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N10
cycloneive_lcell_comb \Mux52~10 (
// Equation(s):
// \Mux52~10_combout  = (dcifimemload_19 & (((\my_reg[25][11]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[17][11]~q  & ((!dcifimemload_18))))

	.dataa(\my_reg[17][11]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[25][11]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux52~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~10 .lut_mask = 16'hCCE2;
defparam \Mux52~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N14
cycloneive_lcell_comb \Mux52~11 (
// Equation(s):
// \Mux52~11_combout  = (\Mux52~10_combout  & ((\my_reg[29][11]~q ) # ((!dcifimemload_18)))) # (!\Mux52~10_combout  & (((\my_reg[21][11]~q  & dcifimemload_18))))

	.dataa(\my_reg[29][11]~q ),
	.datab(\my_reg[21][11]~q ),
	.datac(\Mux52~10_combout ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux52~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~11 .lut_mask = 16'hACF0;
defparam \Mux52~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N20
cycloneive_lcell_comb \Mux52~14 (
// Equation(s):
// \Mux52~14_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[20][11]~q ))) # (!dcifimemload_18 & (\my_reg[16][11]~q ))))

	.dataa(\my_reg[16][11]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[20][11]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux52~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~14 .lut_mask = 16'hFC22;
defparam \Mux52~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N26
cycloneive_lcell_comb \Mux52~15 (
// Equation(s):
// \Mux52~15_combout  = (dcifimemload_19 & ((\Mux52~14_combout  & (\my_reg[28][11]~q )) # (!\Mux52~14_combout  & ((\my_reg[24][11]~q ))))) # (!dcifimemload_19 & (((\Mux52~14_combout ))))

	.dataa(\my_reg[28][11]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[24][11]~q ),
	.datad(\Mux52~14_combout ),
	.cin(gnd),
	.combout(\Mux52~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~15 .lut_mask = 16'hBBC0;
defparam \Mux52~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y42_N11
dffeas \my_reg[26][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][11] .is_wysiwyg = "true";
defparam \my_reg[26][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y42_N1
dffeas \my_reg[22][11] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][11] .is_wysiwyg = "true";
defparam \my_reg[22][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N0
cycloneive_lcell_comb \Mux52~12 (
// Equation(s):
// \Mux52~12_combout  = (dcifimemload_18 & (((\my_reg[22][11]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[18][11]~q  & ((!dcifimemload_19))))

	.dataa(\my_reg[18][11]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[22][11]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux52~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~12 .lut_mask = 16'hCCE2;
defparam \Mux52~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N10
cycloneive_lcell_comb \Mux52~13 (
// Equation(s):
// \Mux52~13_combout  = (dcifimemload_19 & ((\Mux52~12_combout  & (\my_reg[30][11]~q )) # (!\Mux52~12_combout  & ((\my_reg[26][11]~q ))))) # (!dcifimemload_19 & (((\Mux52~12_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[30][11]~q ),
	.datac(\my_reg[26][11]~q ),
	.datad(\Mux52~12_combout ),
	.cin(gnd),
	.combout(\Mux52~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~13 .lut_mask = 16'hDDA0;
defparam \Mux52~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N10
cycloneive_lcell_comb \Mux52~16 (
// Equation(s):
// \Mux52~16_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux52~13_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & (\Mux52~15_combout )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux52~15_combout ),
	.datad(\Mux52~13_combout ),
	.cin(gnd),
	.combout(\Mux52~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~16 .lut_mask = 16'hBA98;
defparam \Mux52~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N15
dffeas \my_reg[23][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][10] .is_wysiwyg = "true";
defparam \my_reg[23][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N4
cycloneive_lcell_comb \my_reg[19][10]~feeder (
// Equation(s):
// \my_reg[19][10]~feeder_combout  = \wdat~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat23),
	.cin(gnd),
	.combout(\my_reg[19][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[19][10]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[19][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N5
dffeas \my_reg[19][10] (
	.clk(CLK),
	.d(\my_reg[19][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][10] .is_wysiwyg = "true";
defparam \my_reg[19][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N2
cycloneive_lcell_comb \Mux21~7 (
// Equation(s):
// \Mux21~7_combout  = (dcifimemload_24 & ((\my_reg[27][10]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\my_reg[19][10]~q  & !dcifimemload_23))))

	.dataa(\my_reg[27][10]~q ),
	.datab(\my_reg[19][10]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux21~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~7 .lut_mask = 16'hF0AC;
defparam \Mux21~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N16
cycloneive_lcell_comb \Mux21~8 (
// Equation(s):
// \Mux21~8_combout  = (dcifimemload_23 & ((\Mux21~7_combout  & (\my_reg[31][10]~q )) # (!\Mux21~7_combout  & ((\my_reg[23][10]~q ))))) # (!dcifimemload_23 & (((\Mux21~7_combout ))))

	.dataa(\my_reg[31][10]~q ),
	.datab(\my_reg[23][10]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux21~7_combout ),
	.cin(gnd),
	.combout(\Mux21~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~8 .lut_mask = 16'hAFC0;
defparam \Mux21~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N13
dffeas \my_reg[29][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][10] .is_wysiwyg = "true";
defparam \my_reg[29][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N15
dffeas \my_reg[21][10] (
	.clk(CLK),
	.d(wdat23),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][10] .is_wysiwyg = "true";
defparam \my_reg[21][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N12
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// \Mux21~1_combout  = (\Mux21~0_combout  & (((\my_reg[29][10]~q )) # (!dcifimemload_23))) # (!\Mux21~0_combout  & (dcifimemload_23 & ((\my_reg[21][10]~q ))))

	.dataa(\Mux21~0_combout ),
	.datab(dcifimemload_23),
	.datac(\my_reg[29][10]~q ),
	.datad(\my_reg[21][10]~q ),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'hE6A2;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N25
dffeas \my_reg[24][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][10] .is_wysiwyg = "true";
defparam \my_reg[24][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N11
dffeas \my_reg[28][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][10] .is_wysiwyg = "true";
defparam \my_reg[28][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y40_N23
dffeas \my_reg[20][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][10] .is_wysiwyg = "true";
defparam \my_reg[20][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N17
dffeas \my_reg[16][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][10] .is_wysiwyg = "true";
defparam \my_reg[16][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N16
cycloneive_lcell_comb \Mux21~4 (
// Equation(s):
// \Mux21~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[20][10]~q )) # (!dcifimemload_23 & ((\my_reg[16][10]~q )))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[20][10]~q ),
	.datac(\my_reg[16][10]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~4 .lut_mask = 16'hEE50;
defparam \Mux21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N10
cycloneive_lcell_comb \Mux21~5 (
// Equation(s):
// \Mux21~5_combout  = (dcifimemload_24 & ((\Mux21~4_combout  & ((\my_reg[28][10]~q ))) # (!\Mux21~4_combout  & (\my_reg[24][10]~q )))) # (!dcifimemload_24 & (((\Mux21~4_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[24][10]~q ),
	.datac(\my_reg[28][10]~q ),
	.datad(\Mux21~4_combout ),
	.cin(gnd),
	.combout(\Mux21~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~5 .lut_mask = 16'hF588;
defparam \Mux21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N29
dffeas \my_reg[30][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][10] .is_wysiwyg = "true";
defparam \my_reg[30][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N25
dffeas \my_reg[18][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][10] .is_wysiwyg = "true";
defparam \my_reg[18][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N24
cycloneive_lcell_comb \Mux21~2 (
// Equation(s):
// \Mux21~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[22][10]~q )) # (!dcifimemload_23 & ((\my_reg[18][10]~q )))))

	.dataa(\my_reg[22][10]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[18][10]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~2 .lut_mask = 16'hEE30;
defparam \Mux21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N28
cycloneive_lcell_comb \Mux21~3 (
// Equation(s):
// \Mux21~3_combout  = (dcifimemload_24 & ((\Mux21~2_combout  & ((\my_reg[30][10]~q ))) # (!\Mux21~2_combout  & (\my_reg[26][10]~q )))) # (!dcifimemload_24 & (((\Mux21~2_combout ))))

	.dataa(\my_reg[26][10]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[30][10]~q ),
	.datad(\Mux21~2_combout ),
	.cin(gnd),
	.combout(\Mux21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~3 .lut_mask = 16'hF388;
defparam \Mux21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N24
cycloneive_lcell_comb \Mux21~6 (
// Equation(s):
// \Mux21~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux21~3_combout ))) # (!dcifimemload_22 & (\Mux21~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux21~5_combout ),
	.datad(\Mux21~3_combout ),
	.cin(gnd),
	.combout(\Mux21~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~6 .lut_mask = 16'hDC98;
defparam \Mux21~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N26
cycloneive_lcell_comb \Mux21~9 (
// Equation(s):
// \Mux21~9_combout  = (dcifimemload_21 & ((\Mux21~6_combout  & (\Mux21~8_combout )) # (!\Mux21~6_combout  & ((\Mux21~1_combout ))))) # (!dcifimemload_21 & (((\Mux21~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux21~8_combout ),
	.datac(\Mux21~1_combout ),
	.datad(\Mux21~6_combout ),
	.cin(gnd),
	.combout(\Mux21~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~9 .lut_mask = 16'hDDA0;
defparam \Mux21~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N7
dffeas \my_reg[7][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][10] .is_wysiwyg = "true";
defparam \my_reg[7][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N13
dffeas \my_reg[6][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][10] .is_wysiwyg = "true";
defparam \my_reg[6][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N25
dffeas \my_reg[4][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][10] .is_wysiwyg = "true";
defparam \my_reg[4][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N11
dffeas \my_reg[5][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][10] .is_wysiwyg = "true";
defparam \my_reg[5][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N10
cycloneive_lcell_comb \Mux21~10 (
// Equation(s):
// \Mux21~10_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\my_reg[5][10]~q ))) # (!dcifimemload_21 & (\my_reg[4][10]~q ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[4][10]~q ),
	.datac(\my_reg[5][10]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux21~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~10 .lut_mask = 16'hFA44;
defparam \Mux21~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N12
cycloneive_lcell_comb \Mux21~11 (
// Equation(s):
// \Mux21~11_combout  = (dcifimemload_22 & ((\Mux21~10_combout  & (\my_reg[7][10]~q )) # (!\Mux21~10_combout  & ((\my_reg[6][10]~q ))))) # (!dcifimemload_22 & (((\Mux21~10_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[7][10]~q ),
	.datac(\my_reg[6][10]~q ),
	.datad(\Mux21~10_combout ),
	.cin(gnd),
	.combout(\Mux21~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~11 .lut_mask = 16'hDDA0;
defparam \Mux21~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N11
dffeas \my_reg[2][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][10] .is_wysiwyg = "true";
defparam \my_reg[2][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N17
dffeas \my_reg[1][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][10] .is_wysiwyg = "true";
defparam \my_reg[1][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N19
dffeas \my_reg[3][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][10] .is_wysiwyg = "true";
defparam \my_reg[3][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N18
cycloneive_lcell_comb \Mux21~14 (
// Equation(s):
// \Mux21~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][10]~q ))) # (!dcifimemload_22 & (\my_reg[1][10]~q ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[1][10]~q ),
	.datac(\my_reg[3][10]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux21~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~14 .lut_mask = 16'hA088;
defparam \Mux21~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N4
cycloneive_lcell_comb \Mux21~15 (
// Equation(s):
// \Mux21~15_combout  = (\Mux21~14_combout ) # ((!dcifimemload_21 & (dcifimemload_22 & \my_reg[2][10]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\my_reg[2][10]~q ),
	.datad(\Mux21~14_combout ),
	.cin(gnd),
	.combout(\Mux21~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~15 .lut_mask = 16'hFF40;
defparam \Mux21~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N24
cycloneive_lcell_comb \my_reg[9][10]~feeder (
// Equation(s):
// \my_reg[9][10]~feeder_combout  = \wdat~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat23),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[9][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[9][10]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[9][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y31_N25
dffeas \my_reg[9][10] (
	.clk(CLK),
	.d(\my_reg[9][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][10] .is_wysiwyg = "true";
defparam \my_reg[9][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N19
dffeas \my_reg[11][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][10] .is_wysiwyg = "true";
defparam \my_reg[11][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N21
dffeas \my_reg[8][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][10] .is_wysiwyg = "true";
defparam \my_reg[8][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N20
cycloneive_lcell_comb \Mux21~12 (
// Equation(s):
// \Mux21~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][10]~q )) # (!dcifimemload_22 & ((\my_reg[8][10]~q )))))

	.dataa(\my_reg[10][10]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[8][10]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux21~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~12 .lut_mask = 16'hEE30;
defparam \Mux21~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N18
cycloneive_lcell_comb \Mux21~13 (
// Equation(s):
// \Mux21~13_combout  = (dcifimemload_21 & ((\Mux21~12_combout  & ((\my_reg[11][10]~q ))) # (!\Mux21~12_combout  & (\my_reg[9][10]~q )))) # (!dcifimemload_21 & (((\Mux21~12_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][10]~q ),
	.datac(\my_reg[11][10]~q ),
	.datad(\Mux21~12_combout ),
	.cin(gnd),
	.combout(\Mux21~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~13 .lut_mask = 16'hF588;
defparam \Mux21~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N22
cycloneive_lcell_comb \Mux21~16 (
// Equation(s):
// \Mux21~16_combout  = (dcifimemload_24 & ((dcifimemload_23) # ((\Mux21~13_combout )))) # (!dcifimemload_24 & (!dcifimemload_23 & (\Mux21~15_combout )))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux21~15_combout ),
	.datad(\Mux21~13_combout ),
	.cin(gnd),
	.combout(\Mux21~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~16 .lut_mask = 16'hBA98;
defparam \Mux21~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N22
cycloneive_lcell_comb \my_reg[15][10]~feeder (
// Equation(s):
// \my_reg[15][10]~feeder_combout  = \wdat~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat23),
	.cin(gnd),
	.combout(\my_reg[15][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[15][10]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[15][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N23
dffeas \my_reg[15][10] (
	.clk(CLK),
	.d(\my_reg[15][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][10] .is_wysiwyg = "true";
defparam \my_reg[15][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N5
dffeas \my_reg[12][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][10] .is_wysiwyg = "true";
defparam \my_reg[12][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N8
cycloneive_lcell_comb \Mux21~17 (
// Equation(s):
// \Mux21~17_combout  = (dcifimemload_21 & ((\my_reg[13][10]~q ) # ((dcifimemload_22)))) # (!dcifimemload_21 & (((\my_reg[12][10]~q  & !dcifimemload_22))))

	.dataa(\my_reg[13][10]~q ),
	.datab(\my_reg[12][10]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux21~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~17 .lut_mask = 16'hF0AC;
defparam \Mux21~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N6
cycloneive_lcell_comb \Mux21~18 (
// Equation(s):
// \Mux21~18_combout  = (\Mux21~17_combout  & (((\my_reg[15][10]~q ) # (!dcifimemload_22)))) # (!\Mux21~17_combout  & (\my_reg[14][10]~q  & ((dcifimemload_22))))

	.dataa(\my_reg[14][10]~q ),
	.datab(\my_reg[15][10]~q ),
	.datac(\Mux21~17_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux21~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~18 .lut_mask = 16'hCAF0;
defparam \Mux21~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N0
cycloneive_lcell_comb \Mux21~19 (
// Equation(s):
// \Mux21~19_combout  = (dcifimemload_23 & ((\Mux21~16_combout  & ((\Mux21~18_combout ))) # (!\Mux21~16_combout  & (\Mux21~11_combout )))) # (!dcifimemload_23 & (((\Mux21~16_combout ))))

	.dataa(\Mux21~11_combout ),
	.datab(dcifimemload_23),
	.datac(\Mux21~16_combout ),
	.datad(\Mux21~18_combout ),
	.cin(gnd),
	.combout(\Mux21~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~19 .lut_mask = 16'hF838;
defparam \Mux21~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N24
cycloneive_lcell_comb \my_reg[10][10]~feeder (
// Equation(s):
// \my_reg[10][10]~feeder_combout  = \wdat~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat23),
	.cin(gnd),
	.combout(\my_reg[10][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[10][10]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[10][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y31_N25
dffeas \my_reg[10][10] (
	.clk(CLK),
	.d(\my_reg[10][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][10] .is_wysiwyg = "true";
defparam \my_reg[10][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N10
cycloneive_lcell_comb \Mux53~0 (
// Equation(s):
// \Mux53~0_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[10][10]~q ))) # (!dcifimemload_17 & (\my_reg[8][10]~q ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[8][10]~q ),
	.datac(\my_reg[10][10]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux53~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~0 .lut_mask = 16'hFA44;
defparam \Mux53~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N8
cycloneive_lcell_comb \Mux53~1 (
// Equation(s):
// \Mux53~1_combout  = (dcifimemload_16 & ((\Mux53~0_combout  & (\my_reg[11][10]~q )) # (!\Mux53~0_combout  & ((\my_reg[9][10]~q ))))) # (!dcifimemload_16 & (((\Mux53~0_combout ))))

	.dataa(\my_reg[11][10]~q ),
	.datab(\my_reg[9][10]~q ),
	.datac(dcifimemload_16),
	.datad(\Mux53~0_combout ),
	.cin(gnd),
	.combout(\Mux53~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~1 .lut_mask = 16'hAFC0;
defparam \Mux53~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N16
cycloneive_lcell_comb \Mux53~4 (
// Equation(s):
// \Mux53~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\my_reg[3][10]~q )) # (!dcifimemload_17 & ((\my_reg[1][10]~q )))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[3][10]~q ),
	.datac(\my_reg[1][10]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux53~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~4 .lut_mask = 16'hD800;
defparam \Mux53~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N10
cycloneive_lcell_comb \Mux53~5 (
// Equation(s):
// \Mux53~5_combout  = (\Mux53~4_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \my_reg[2][10]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\my_reg[2][10]~q ),
	.datad(\Mux53~4_combout ),
	.cin(gnd),
	.combout(\Mux53~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~5 .lut_mask = 16'hFF20;
defparam \Mux53~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N24
cycloneive_lcell_comb \Mux53~2 (
// Equation(s):
// \Mux53~2_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\my_reg[5][10]~q )) # (!dcifimemload_16 & ((\my_reg[4][10]~q )))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[5][10]~q ),
	.datac(\my_reg[4][10]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux53~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~2 .lut_mask = 16'hEE50;
defparam \Mux53~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N6
cycloneive_lcell_comb \Mux53~3 (
// Equation(s):
// \Mux53~3_combout  = (\Mux53~2_combout  & (((\my_reg[7][10]~q ) # (!dcifimemload_17)))) # (!\Mux53~2_combout  & (\my_reg[6][10]~q  & ((dcifimemload_17))))

	.dataa(\my_reg[6][10]~q ),
	.datab(\Mux53~2_combout ),
	.datac(\my_reg[7][10]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux53~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~3 .lut_mask = 16'hE2CC;
defparam \Mux53~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N30
cycloneive_lcell_comb \Mux53~6 (
// Equation(s):
// \Mux53~6_combout  = (dcifimemload_18 & ((dcifimemload_19) # ((\Mux53~3_combout )))) # (!dcifimemload_18 & (!dcifimemload_19 & (\Mux53~5_combout )))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux53~5_combout ),
	.datad(\Mux53~3_combout ),
	.cin(gnd),
	.combout(\Mux53~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~6 .lut_mask = 16'hBA98;
defparam \Mux53~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N12
cycloneive_lcell_comb \my_reg[14][10]~feeder (
// Equation(s):
// \my_reg[14][10]~feeder_combout  = \wdat~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat23),
	.cin(gnd),
	.combout(\my_reg[14][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[14][10]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[14][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N13
dffeas \my_reg[14][10] (
	.clk(CLK),
	.d(\my_reg[14][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][10] .is_wysiwyg = "true";
defparam \my_reg[14][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N14
cycloneive_lcell_comb \my_reg[13][10]~feeder (
// Equation(s):
// \my_reg[13][10]~feeder_combout  = \wdat~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat23),
	.cin(gnd),
	.combout(\my_reg[13][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[13][10]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[13][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N15
dffeas \my_reg[13][10] (
	.clk(CLK),
	.d(\my_reg[13][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][10] .is_wysiwyg = "true";
defparam \my_reg[13][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N4
cycloneive_lcell_comb \Mux53~7 (
// Equation(s):
// \Mux53~7_combout  = (dcifimemload_17 & (dcifimemload_16)) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[13][10]~q ))) # (!dcifimemload_16 & (\my_reg[12][10]~q ))))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\my_reg[12][10]~q ),
	.datad(\my_reg[13][10]~q ),
	.cin(gnd),
	.combout(\Mux53~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~7 .lut_mask = 16'hDC98;
defparam \Mux53~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N16
cycloneive_lcell_comb \Mux53~8 (
// Equation(s):
// \Mux53~8_combout  = (\Mux53~7_combout  & (((\my_reg[15][10]~q ) # (!dcifimemload_17)))) # (!\Mux53~7_combout  & (\my_reg[14][10]~q  & ((dcifimemload_17))))

	.dataa(\my_reg[14][10]~q ),
	.datab(\my_reg[15][10]~q ),
	.datac(\Mux53~7_combout ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux53~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~8 .lut_mask = 16'hCAF0;
defparam \Mux53~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N23
dffeas \my_reg[25][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][10] .is_wysiwyg = "true";
defparam \my_reg[25][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N18
cycloneive_lcell_comb \Mux53~10 (
// Equation(s):
// \Mux53~10_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[21][10]~q ))) # (!dcifimemload_18 & (\my_reg[17][10]~q ))))

	.dataa(\my_reg[17][10]~q ),
	.datab(\my_reg[21][10]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux53~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~10 .lut_mask = 16'hFC0A;
defparam \Mux53~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N22
cycloneive_lcell_comb \Mux53~11 (
// Equation(s):
// \Mux53~11_combout  = (dcifimemload_19 & ((\Mux53~10_combout  & (\my_reg[29][10]~q )) # (!\Mux53~10_combout  & ((\my_reg[25][10]~q ))))) # (!dcifimemload_19 & (((\Mux53~10_combout ))))

	.dataa(\my_reg[29][10]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[25][10]~q ),
	.datad(\Mux53~10_combout ),
	.cin(gnd),
	.combout(\Mux53~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~11 .lut_mask = 16'hBBC0;
defparam \Mux53~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N24
cycloneive_lcell_comb \my_reg[31][10]~feeder (
// Equation(s):
// \my_reg[31][10]~feeder_combout  = \wdat~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat23),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[31][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[31][10]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[31][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N25
dffeas \my_reg[31][10] (
	.clk(CLK),
	.d(\my_reg[31][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][10] .is_wysiwyg = "true";
defparam \my_reg[31][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y36_N23
dffeas \my_reg[27][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][10] .is_wysiwyg = "true";
defparam \my_reg[27][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N14
cycloneive_lcell_comb \Mux53~17 (
// Equation(s):
// \Mux53~17_combout  = (dcifimemload_19 & (dcifimemload_18)) # (!dcifimemload_19 & ((dcifimemload_18 & (\my_reg[23][10]~q )) # (!dcifimemload_18 & ((\my_reg[19][10]~q )))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\my_reg[23][10]~q ),
	.datad(\my_reg[19][10]~q ),
	.cin(gnd),
	.combout(\Mux53~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~17 .lut_mask = 16'hD9C8;
defparam \Mux53~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N22
cycloneive_lcell_comb \Mux53~18 (
// Equation(s):
// \Mux53~18_combout  = (dcifimemload_19 & ((\Mux53~17_combout  & (\my_reg[31][10]~q )) # (!\Mux53~17_combout  & ((\my_reg[27][10]~q ))))) # (!dcifimemload_19 & (((\Mux53~17_combout ))))

	.dataa(\my_reg[31][10]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[27][10]~q ),
	.datad(\Mux53~17_combout ),
	.cin(gnd),
	.combout(\Mux53~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~18 .lut_mask = 16'hBBC0;
defparam \Mux53~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N24
cycloneive_lcell_comb \Mux53~14 (
// Equation(s):
// \Mux53~14_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[24][10]~q ))) # (!dcifimemload_19 & (\my_reg[16][10]~q ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[16][10]~q ),
	.datac(\my_reg[24][10]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux53~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~14 .lut_mask = 16'hFA44;
defparam \Mux53~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N22
cycloneive_lcell_comb \Mux53~15 (
// Equation(s):
// \Mux53~15_combout  = (dcifimemload_18 & ((\Mux53~14_combout  & (\my_reg[28][10]~q )) # (!\Mux53~14_combout  & ((\my_reg[20][10]~q ))))) # (!dcifimemload_18 & (((\Mux53~14_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[28][10]~q ),
	.datac(\my_reg[20][10]~q ),
	.datad(\Mux53~14_combout ),
	.cin(gnd),
	.combout(\Mux53~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~15 .lut_mask = 16'hDDA0;
defparam \Mux53~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N3
dffeas \my_reg[22][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][10] .is_wysiwyg = "true";
defparam \my_reg[22][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N23
dffeas \my_reg[26][10] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][10] .is_wysiwyg = "true";
defparam \my_reg[26][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N22
cycloneive_lcell_comb \Mux53~12 (
// Equation(s):
// \Mux53~12_combout  = (dcifimemload_19 & (((\my_reg[26][10]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[18][10]~q  & ((!dcifimemload_18))))

	.dataa(\my_reg[18][10]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[26][10]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux53~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~12 .lut_mask = 16'hCCE2;
defparam \Mux53~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N2
cycloneive_lcell_comb \Mux53~13 (
// Equation(s):
// \Mux53~13_combout  = (dcifimemload_18 & ((\Mux53~12_combout  & (\my_reg[30][10]~q )) # (!\Mux53~12_combout  & ((\my_reg[22][10]~q ))))) # (!dcifimemload_18 & (((\Mux53~12_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[30][10]~q ),
	.datac(\my_reg[22][10]~q ),
	.datad(\Mux53~12_combout ),
	.cin(gnd),
	.combout(\Mux53~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~13 .lut_mask = 16'hDDA0;
defparam \Mux53~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N20
cycloneive_lcell_comb \Mux53~16 (
// Equation(s):
// \Mux53~16_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux53~13_combout ))) # (!dcifimemload_17 & (\Mux53~15_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux53~15_combout ),
	.datad(\Mux53~13_combout ),
	.cin(gnd),
	.combout(\Mux53~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~16 .lut_mask = 16'hDC98;
defparam \Mux53~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N29
dffeas \my_reg[25][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][9] .is_wysiwyg = "true";
defparam \my_reg[25][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N9
dffeas \my_reg[29][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][9] .is_wysiwyg = "true";
defparam \my_reg[29][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N8
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// \Mux22~1_combout  = (\Mux22~0_combout  & (((\my_reg[29][9]~q ) # (!dcifimemload_24)))) # (!\Mux22~0_combout  & (\my_reg[25][9]~q  & ((dcifimemload_24))))

	.dataa(\Mux22~0_combout ),
	.datab(\my_reg[25][9]~q ),
	.datac(\my_reg[29][9]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'hE4AA;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N4
cycloneive_lcell_comb \my_reg[27][9]~feeder (
// Equation(s):
// \my_reg[27][9]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat24),
	.cin(gnd),
	.combout(\my_reg[27][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[27][9]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[27][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N5
dffeas \my_reg[27][9] (
	.clk(CLK),
	.d(\my_reg[27][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][9] .is_wysiwyg = "true";
defparam \my_reg[27][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N31
dffeas \my_reg[31][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][9] .is_wysiwyg = "true";
defparam \my_reg[31][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N14
cycloneive_lcell_comb \my_reg[19][9]~feeder (
// Equation(s):
// \my_reg[19][9]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat24),
	.cin(gnd),
	.combout(\my_reg[19][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[19][9]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[19][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N15
dffeas \my_reg[19][9] (
	.clk(CLK),
	.d(\my_reg[19][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][9] .is_wysiwyg = "true";
defparam \my_reg[19][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N29
dffeas \my_reg[23][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][9] .is_wysiwyg = "true";
defparam \my_reg[23][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N28
cycloneive_lcell_comb \Mux22~7 (
// Equation(s):
// \Mux22~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\my_reg[23][9]~q ))) # (!dcifimemload_23 & (\my_reg[19][9]~q ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[19][9]~q ),
	.datac(\my_reg[23][9]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux22~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~7 .lut_mask = 16'hFA44;
defparam \Mux22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N30
cycloneive_lcell_comb \Mux22~8 (
// Equation(s):
// \Mux22~8_combout  = (dcifimemload_24 & ((\Mux22~7_combout  & ((\my_reg[31][9]~q ))) # (!\Mux22~7_combout  & (\my_reg[27][9]~q )))) # (!dcifimemload_24 & (((\Mux22~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[27][9]~q ),
	.datac(\my_reg[31][9]~q ),
	.datad(\Mux22~7_combout ),
	.cin(gnd),
	.combout(\Mux22~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~8 .lut_mask = 16'hF588;
defparam \Mux22~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N8
cycloneive_lcell_comb \my_reg[28][9]~feeder (
// Equation(s):
// \my_reg[28][9]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat24),
	.cin(gnd),
	.combout(\my_reg[28][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[28][9]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[28][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N9
dffeas \my_reg[28][9] (
	.clk(CLK),
	.d(\my_reg[28][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][9] .is_wysiwyg = "true";
defparam \my_reg[28][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N28
cycloneive_lcell_comb \my_reg[16][9]~feeder (
// Equation(s):
// \my_reg[16][9]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat24),
	.cin(gnd),
	.combout(\my_reg[16][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[16][9]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[16][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N29
dffeas \my_reg[16][9] (
	.clk(CLK),
	.d(\my_reg[16][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][9] .is_wysiwyg = "true";
defparam \my_reg[16][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N22
cycloneive_lcell_comb \Mux22~4 (
// Equation(s):
// \Mux22~4_combout  = (dcifimemload_24 & ((\my_reg[24][9]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\my_reg[16][9]~q  & !dcifimemload_23))))

	.dataa(\my_reg[24][9]~q ),
	.datab(\my_reg[16][9]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~4 .lut_mask = 16'hF0AC;
defparam \Mux22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N14
cycloneive_lcell_comb \Mux22~5 (
// Equation(s):
// \Mux22~5_combout  = (\Mux22~4_combout  & (((\my_reg[28][9]~q ) # (!dcifimemload_23)))) # (!\Mux22~4_combout  & (\my_reg[20][9]~q  & ((dcifimemload_23))))

	.dataa(\my_reg[20][9]~q ),
	.datab(\my_reg[28][9]~q ),
	.datac(\Mux22~4_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux22~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~5 .lut_mask = 16'hCAF0;
defparam \Mux22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y42_N17
dffeas \my_reg[22][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][9] .is_wysiwyg = "true";
defparam \my_reg[22][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N16
cycloneive_lcell_comb \my_reg[18][9]~feeder (
// Equation(s):
// \my_reg[18][9]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat24),
	.cin(gnd),
	.combout(\my_reg[18][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[18][9]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[18][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N17
dffeas \my_reg[18][9] (
	.clk(CLK),
	.d(\my_reg[18][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][9] .is_wysiwyg = "true";
defparam \my_reg[18][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N6
cycloneive_lcell_comb \Mux22~2 (
// Equation(s):
// \Mux22~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[26][9]~q )) # (!dcifimemload_24 & ((\my_reg[18][9]~q )))))

	.dataa(\my_reg[26][9]~q ),
	.datab(\my_reg[18][9]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~2 .lut_mask = 16'hFA0C;
defparam \Mux22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N2
cycloneive_lcell_comb \Mux22~3 (
// Equation(s):
// \Mux22~3_combout  = (dcifimemload_23 & ((\Mux22~2_combout  & (\my_reg[30][9]~q )) # (!\Mux22~2_combout  & ((\my_reg[22][9]~q ))))) # (!dcifimemload_23 & (((\Mux22~2_combout ))))

	.dataa(\my_reg[30][9]~q ),
	.datab(\my_reg[22][9]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux22~2_combout ),
	.cin(gnd),
	.combout(\Mux22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~3 .lut_mask = 16'hAFC0;
defparam \Mux22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N28
cycloneive_lcell_comb \Mux22~6 (
// Equation(s):
// \Mux22~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux22~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & (\Mux22~5_combout )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux22~5_combout ),
	.datad(\Mux22~3_combout ),
	.cin(gnd),
	.combout(\Mux22~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~6 .lut_mask = 16'hBA98;
defparam \Mux22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N14
cycloneive_lcell_comb \Mux22~9 (
// Equation(s):
// \Mux22~9_combout  = (dcifimemload_21 & ((\Mux22~6_combout  & ((\Mux22~8_combout ))) # (!\Mux22~6_combout  & (\Mux22~1_combout )))) # (!dcifimemload_21 & (((\Mux22~6_combout ))))

	.dataa(\Mux22~1_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux22~8_combout ),
	.datad(\Mux22~6_combout ),
	.cin(gnd),
	.combout(\Mux22~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~9 .lut_mask = 16'hF388;
defparam \Mux22~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N27
dffeas \my_reg[14][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][9] .is_wysiwyg = "true";
defparam \my_reg[14][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N1
dffeas \my_reg[13][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][9] .is_wysiwyg = "true";
defparam \my_reg[13][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N0
cycloneive_lcell_comb \Mux22~17 (
// Equation(s):
// \Mux22~17_combout  = (dcifimemload_21 & (((\my_reg[13][9]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\my_reg[12][9]~q  & ((!dcifimemload_22))))

	.dataa(\my_reg[12][9]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[13][9]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux22~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~17 .lut_mask = 16'hCCE2;
defparam \Mux22~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N10
cycloneive_lcell_comb \Mux22~18 (
// Equation(s):
// \Mux22~18_combout  = (dcifimemload_22 & ((\Mux22~17_combout  & (\my_reg[15][9]~q )) # (!\Mux22~17_combout  & ((\my_reg[14][9]~q ))))) # (!dcifimemload_22 & (((\Mux22~17_combout ))))

	.dataa(\my_reg[15][9]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[14][9]~q ),
	.datad(\Mux22~17_combout ),
	.cin(gnd),
	.combout(\Mux22~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~18 .lut_mask = 16'hBBC0;
defparam \Mux22~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N31
dffeas \my_reg[11][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][9] .is_wysiwyg = "true";
defparam \my_reg[11][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N9
dffeas \my_reg[8][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][9] .is_wysiwyg = "true";
defparam \my_reg[8][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N19
dffeas \my_reg[10][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][9] .is_wysiwyg = "true";
defparam \my_reg[10][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N18
cycloneive_lcell_comb \Mux22~10 (
// Equation(s):
// \Mux22~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[10][9]~q ))) # (!dcifimemload_22 & (\my_reg[8][9]~q ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[8][9]~q ),
	.datac(\my_reg[10][9]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux22~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~10 .lut_mask = 16'hFA44;
defparam \Mux22~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N20
cycloneive_lcell_comb \Mux22~11 (
// Equation(s):
// \Mux22~11_combout  = (dcifimemload_21 & ((\Mux22~10_combout  & ((\my_reg[11][9]~q ))) # (!\Mux22~10_combout  & (\my_reg[9][9]~q )))) # (!dcifimemload_21 & (((\Mux22~10_combout ))))

	.dataa(\my_reg[9][9]~q ),
	.datab(\my_reg[11][9]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux22~10_combout ),
	.cin(gnd),
	.combout(\Mux22~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~11 .lut_mask = 16'hCFA0;
defparam \Mux22~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y32_N25
dffeas \my_reg[6][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][9] .is_wysiwyg = "true";
defparam \my_reg[6][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N3
dffeas \my_reg[7][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][9] .is_wysiwyg = "true";
defparam \my_reg[7][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N25
dffeas \my_reg[4][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][9] .is_wysiwyg = "true";
defparam \my_reg[4][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N24
cycloneive_lcell_comb \Mux22~12 (
// Equation(s):
// \Mux22~12_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\my_reg[5][9]~q )) # (!dcifimemload_21 & ((\my_reg[4][9]~q )))))

	.dataa(\my_reg[5][9]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[4][9]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux22~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~12 .lut_mask = 16'hEE30;
defparam \Mux22~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N2
cycloneive_lcell_comb \Mux22~13 (
// Equation(s):
// \Mux22~13_combout  = (dcifimemload_22 & ((\Mux22~12_combout  & ((\my_reg[7][9]~q ))) # (!\Mux22~12_combout  & (\my_reg[6][9]~q )))) # (!dcifimemload_22 & (((\Mux22~12_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[6][9]~q ),
	.datac(\my_reg[7][9]~q ),
	.datad(\Mux22~12_combout ),
	.cin(gnd),
	.combout(\Mux22~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~13 .lut_mask = 16'hF588;
defparam \Mux22~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N13
dffeas \my_reg[1][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][9] .is_wysiwyg = "true";
defparam \my_reg[1][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N17
dffeas \my_reg[3][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][9] .is_wysiwyg = "true";
defparam \my_reg[3][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N16
cycloneive_lcell_comb \Mux22~14 (
// Equation(s):
// \Mux22~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][9]~q ))) # (!dcifimemload_22 & (\my_reg[1][9]~q ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[1][9]~q ),
	.datac(\my_reg[3][9]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux22~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~14 .lut_mask = 16'hA088;
defparam \Mux22~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N28
cycloneive_lcell_comb \Mux22~15 (
// Equation(s):
// \Mux22~15_combout  = (\Mux22~14_combout ) # ((\my_reg[2][9]~q  & (dcifimemload_22 & !dcifimemload_21)))

	.dataa(\my_reg[2][9]~q ),
	.datab(dcifimemload_22),
	.datac(dcifimemload_21),
	.datad(\Mux22~14_combout ),
	.cin(gnd),
	.combout(\Mux22~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~15 .lut_mask = 16'hFF08;
defparam \Mux22~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N2
cycloneive_lcell_comb \Mux22~16 (
// Equation(s):
// \Mux22~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & (\Mux22~13_combout )) # (!dcifimemload_23 & ((\Mux22~15_combout )))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux22~13_combout ),
	.datad(\Mux22~15_combout ),
	.cin(gnd),
	.combout(\Mux22~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~16 .lut_mask = 16'hD9C8;
defparam \Mux22~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N20
cycloneive_lcell_comb \Mux22~19 (
// Equation(s):
// \Mux22~19_combout  = (dcifimemload_24 & ((\Mux22~16_combout  & (\Mux22~18_combout )) # (!\Mux22~16_combout  & ((\Mux22~11_combout ))))) # (!dcifimemload_24 & (((\Mux22~16_combout ))))

	.dataa(\Mux22~18_combout ),
	.datab(\Mux22~11_combout ),
	.datac(dcifimemload_24),
	.datad(\Mux22~16_combout ),
	.cin(gnd),
	.combout(\Mux22~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~19 .lut_mask = 16'hAFC0;
defparam \Mux22~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N8
cycloneive_lcell_comb \Mux54~2 (
// Equation(s):
// \Mux54~2_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\my_reg[10][9]~q )) # (!dcifimemload_17 & ((\my_reg[8][9]~q )))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[10][9]~q ),
	.datac(\my_reg[8][9]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux54~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~2 .lut_mask = 16'hEE50;
defparam \Mux54~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N30
cycloneive_lcell_comb \Mux54~3 (
// Equation(s):
// \Mux54~3_combout  = (\Mux54~2_combout  & (((\my_reg[11][9]~q ) # (!dcifimemload_16)))) # (!\Mux54~2_combout  & (\my_reg[9][9]~q  & ((dcifimemload_16))))

	.dataa(\my_reg[9][9]~q ),
	.datab(\Mux54~2_combout ),
	.datac(\my_reg[11][9]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux54~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~3 .lut_mask = 16'hE2CC;
defparam \Mux54~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y33_N9
dffeas \my_reg[2][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][9] .is_wysiwyg = "true";
defparam \my_reg[2][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N12
cycloneive_lcell_comb \Mux54~4 (
// Equation(s):
// \Mux54~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\my_reg[3][9]~q )) # (!dcifimemload_17 & ((\my_reg[1][9]~q )))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[3][9]~q ),
	.datac(\my_reg[1][9]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux54~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~4 .lut_mask = 16'hD800;
defparam \Mux54~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N8
cycloneive_lcell_comb \Mux54~5 (
// Equation(s):
// \Mux54~5_combout  = (\Mux54~4_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \my_reg[2][9]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\my_reg[2][9]~q ),
	.datad(\Mux54~4_combout ),
	.cin(gnd),
	.combout(\Mux54~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~5 .lut_mask = 16'hFF20;
defparam \Mux54~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N10
cycloneive_lcell_comb \Mux54~6 (
// Equation(s):
// \Mux54~6_combout  = (dcifimemload_19 & ((\Mux54~3_combout ) # ((dcifimemload_18)))) # (!dcifimemload_19 & (((\Mux54~5_combout  & !dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\Mux54~3_combout ),
	.datac(\Mux54~5_combout ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux54~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~6 .lut_mask = 16'hAAD8;
defparam \Mux54~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N30
cycloneive_lcell_comb \my_reg[15][9]~feeder (
// Equation(s):
// \my_reg[15][9]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat24),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[15][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[15][9]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[15][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y41_N31
dffeas \my_reg[15][9] (
	.clk(CLK),
	.d(\my_reg[15][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][9] .is_wysiwyg = "true";
defparam \my_reg[15][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N12
cycloneive_lcell_comb \my_reg[12][9]~feeder (
// Equation(s):
// \my_reg[12][9]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat24),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[12][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[12][9]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[12][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y41_N13
dffeas \my_reg[12][9] (
	.clk(CLK),
	.d(\my_reg[12][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][9] .is_wysiwyg = "true";
defparam \my_reg[12][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N0
cycloneive_lcell_comb \Mux54~7 (
// Equation(s):
// \Mux54~7_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\my_reg[13][9]~q )) # (!dcifimemload_16 & ((\my_reg[12][9]~q )))))

	.dataa(\my_reg[13][9]~q ),
	.datab(\my_reg[12][9]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux54~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~7 .lut_mask = 16'hFA0C;
defparam \Mux54~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N10
cycloneive_lcell_comb \Mux54~8 (
// Equation(s):
// \Mux54~8_combout  = (dcifimemload_17 & ((\Mux54~7_combout  & (\my_reg[15][9]~q )) # (!\Mux54~7_combout  & ((\my_reg[14][9]~q ))))) # (!dcifimemload_17 & (((\Mux54~7_combout ))))

	.dataa(\my_reg[15][9]~q ),
	.datab(\my_reg[14][9]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux54~7_combout ),
	.cin(gnd),
	.combout(\Mux54~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~8 .lut_mask = 16'hAFC0;
defparam \Mux54~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y32_N31
dffeas \my_reg[5][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][9] .is_wysiwyg = "true";
defparam \my_reg[5][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N30
cycloneive_lcell_comb \Mux54~0 (
// Equation(s):
// \Mux54~0_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][9]~q ))) # (!dcifimemload_16 & (\my_reg[4][9]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[4][9]~q ),
	.datac(\my_reg[5][9]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux54~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~0 .lut_mask = 16'hFA44;
defparam \Mux54~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N24
cycloneive_lcell_comb \Mux54~1 (
// Equation(s):
// \Mux54~1_combout  = (\Mux54~0_combout  & ((\my_reg[7][9]~q ) # ((!dcifimemload_17)))) # (!\Mux54~0_combout  & (((\my_reg[6][9]~q  & dcifimemload_17))))

	.dataa(\Mux54~0_combout ),
	.datab(\my_reg[7][9]~q ),
	.datac(\my_reg[6][9]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux54~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~1 .lut_mask = 16'hD8AA;
defparam \Mux54~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N12
cycloneive_lcell_comb \my_reg[21][9]~feeder (
// Equation(s):
// \my_reg[21][9]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat24),
	.cin(gnd),
	.combout(\my_reg[21][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][9]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[21][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y33_N13
dffeas \my_reg[21][9] (
	.clk(CLK),
	.d(\my_reg[21][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][9] .is_wysiwyg = "true";
defparam \my_reg[21][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N28
cycloneive_lcell_comb \Mux54~10 (
// Equation(s):
// \Mux54~10_combout  = (dcifimemload_19 & (((\my_reg[25][9]~q ) # (dcifimemload_18)))) # (!dcifimemload_19 & (\my_reg[17][9]~q  & ((!dcifimemload_18))))

	.dataa(\my_reg[17][9]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[25][9]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux54~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~10 .lut_mask = 16'hCCE2;
defparam \Mux54~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N10
cycloneive_lcell_comb \Mux54~11 (
// Equation(s):
// \Mux54~11_combout  = (dcifimemload_18 & ((\Mux54~10_combout  & ((\my_reg[29][9]~q ))) # (!\Mux54~10_combout  & (\my_reg[21][9]~q )))) # (!dcifimemload_18 & (((\Mux54~10_combout ))))

	.dataa(\my_reg[21][9]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[29][9]~q ),
	.datad(\Mux54~10_combout ),
	.cin(gnd),
	.combout(\Mux54~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~11 .lut_mask = 16'hF388;
defparam \Mux54~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N14
cycloneive_lcell_comb \Mux54~17 (
// Equation(s):
// \Mux54~17_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[27][9]~q ))) # (!dcifimemload_19 & (\my_reg[19][9]~q ))))

	.dataa(\my_reg[19][9]~q ),
	.datab(dcifimemload_18),
	.datac(dcifimemload_19),
	.datad(\my_reg[27][9]~q ),
	.cin(gnd),
	.combout(\Mux54~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~17 .lut_mask = 16'hF2C2;
defparam \Mux54~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N16
cycloneive_lcell_comb \Mux54~18 (
// Equation(s):
// \Mux54~18_combout  = (dcifimemload_18 & ((\Mux54~17_combout  & (\my_reg[31][9]~q )) # (!\Mux54~17_combout  & ((\my_reg[23][9]~q ))))) # (!dcifimemload_18 & (((\Mux54~17_combout ))))

	.dataa(\my_reg[31][9]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[23][9]~q ),
	.datad(\Mux54~17_combout ),
	.cin(gnd),
	.combout(\Mux54~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~18 .lut_mask = 16'hBBC0;
defparam \Mux54~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y42_N3
dffeas \my_reg[26][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][9] .is_wysiwyg = "true";
defparam \my_reg[26][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N16
cycloneive_lcell_comb \Mux54~12 (
// Equation(s):
// \Mux54~12_combout  = (dcifimemload_18 & (((\my_reg[22][9]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[18][9]~q  & ((!dcifimemload_19))))

	.dataa(\my_reg[18][9]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[22][9]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux54~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~12 .lut_mask = 16'hCCE2;
defparam \Mux54~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y42_N2
cycloneive_lcell_comb \Mux54~13 (
// Equation(s):
// \Mux54~13_combout  = (dcifimemload_19 & ((\Mux54~12_combout  & (\my_reg[30][9]~q )) # (!\Mux54~12_combout  & ((\my_reg[26][9]~q ))))) # (!dcifimemload_19 & (((\Mux54~12_combout ))))

	.dataa(\my_reg[30][9]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[26][9]~q ),
	.datad(\Mux54~12_combout ),
	.cin(gnd),
	.combout(\Mux54~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~13 .lut_mask = 16'hBBC0;
defparam \Mux54~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N0
cycloneive_lcell_comb \my_reg[24][9]~feeder (
// Equation(s):
// \my_reg[24][9]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat24),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[24][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[24][9]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[24][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y42_N1
dffeas \my_reg[24][9] (
	.clk(CLK),
	.d(\my_reg[24][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][9] .is_wysiwyg = "true";
defparam \my_reg[24][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y42_N7
dffeas \my_reg[20][9] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][9] .is_wysiwyg = "true";
defparam \my_reg[20][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N6
cycloneive_lcell_comb \Mux54~14 (
// Equation(s):
// \Mux54~14_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[20][9]~q ))) # (!dcifimemload_18 & (\my_reg[16][9]~q ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[16][9]~q ),
	.datac(\my_reg[20][9]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux54~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~14 .lut_mask = 16'hFA44;
defparam \Mux54~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N18
cycloneive_lcell_comb \Mux54~15 (
// Equation(s):
// \Mux54~15_combout  = (dcifimemload_19 & ((\Mux54~14_combout  & ((\my_reg[28][9]~q ))) # (!\Mux54~14_combout  & (\my_reg[24][9]~q )))) # (!dcifimemload_19 & (((\Mux54~14_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[24][9]~q ),
	.datac(\my_reg[28][9]~q ),
	.datad(\Mux54~14_combout ),
	.cin(gnd),
	.combout(\Mux54~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~15 .lut_mask = 16'hF588;
defparam \Mux54~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N20
cycloneive_lcell_comb \Mux54~16 (
// Equation(s):
// \Mux54~16_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux54~13_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & ((\Mux54~15_combout ))))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux54~13_combout ),
	.datad(\Mux54~15_combout ),
	.cin(gnd),
	.combout(\Mux54~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~16 .lut_mask = 16'hB9A8;
defparam \Mux54~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N15
dffeas \my_reg[31][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][8] .is_wysiwyg = "true";
defparam \my_reg[31][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N26
cycloneive_lcell_comb \my_reg[19][8]~feeder (
// Equation(s):
// \my_reg[19][8]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat25),
	.cin(gnd),
	.combout(\my_reg[19][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[19][8]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[19][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N27
dffeas \my_reg[19][8] (
	.clk(CLK),
	.d(\my_reg[19][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][8] .is_wysiwyg = "true";
defparam \my_reg[19][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N28
cycloneive_lcell_comb \Mux23~7 (
// Equation(s):
// \Mux23~7_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[27][8]~q )) # (!dcifimemload_24 & ((\my_reg[19][8]~q )))))

	.dataa(\my_reg[27][8]~q ),
	.datab(\my_reg[19][8]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux23~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~7 .lut_mask = 16'hFA0C;
defparam \Mux23~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N14
cycloneive_lcell_comb \Mux23~8 (
// Equation(s):
// \Mux23~8_combout  = (dcifimemload_23 & ((\Mux23~7_combout  & ((\my_reg[31][8]~q ))) # (!\Mux23~7_combout  & (\my_reg[23][8]~q )))) # (!dcifimemload_23 & (((\Mux23~7_combout ))))

	.dataa(\my_reg[23][8]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[31][8]~q ),
	.datad(\Mux23~7_combout ),
	.cin(gnd),
	.combout(\Mux23~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~8 .lut_mask = 16'hF388;
defparam \Mux23~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N31
dffeas \my_reg[29][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][8] .is_wysiwyg = "true";
defparam \my_reg[29][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N19
dffeas \my_reg[25][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][8] .is_wysiwyg = "true";
defparam \my_reg[25][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N16
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (dcifimemload_24 & (((\my_reg[25][8]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\my_reg[17][8]~q  & ((!dcifimemload_23))))

	.dataa(\my_reg[17][8]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[25][8]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hCCE2;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N30
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// \Mux23~1_combout  = (dcifimemload_23 & ((\Mux23~0_combout  & ((\my_reg[29][8]~q ))) # (!\Mux23~0_combout  & (\my_reg[21][8]~q )))) # (!dcifimemload_23 & (((\Mux23~0_combout ))))

	.dataa(\my_reg[21][8]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[29][8]~q ),
	.datad(\Mux23~0_combout ),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'hF388;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N24
cycloneive_lcell_comb \my_reg[30][8]~feeder (
// Equation(s):
// \my_reg[30][8]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat25),
	.cin(gnd),
	.combout(\my_reg[30][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[30][8]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[30][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N25
dffeas \my_reg[30][8] (
	.clk(CLK),
	.d(\my_reg[30][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][8] .is_wysiwyg = "true";
defparam \my_reg[30][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N0
cycloneive_lcell_comb \my_reg[18][8]~feeder (
// Equation(s):
// \my_reg[18][8]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat25),
	.cin(gnd),
	.combout(\my_reg[18][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[18][8]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[18][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N1
dffeas \my_reg[18][8] (
	.clk(CLK),
	.d(\my_reg[18][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][8] .is_wysiwyg = "true";
defparam \my_reg[18][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N18
cycloneive_lcell_comb \Mux23~2 (
// Equation(s):
// \Mux23~2_combout  = (dcifimemload_23 & ((\my_reg[22][8]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[18][8]~q  & !dcifimemload_24))))

	.dataa(\my_reg[22][8]~q ),
	.datab(\my_reg[18][8]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~2 .lut_mask = 16'hF0AC;
defparam \Mux23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N22
cycloneive_lcell_comb \Mux23~3 (
// Equation(s):
// \Mux23~3_combout  = (dcifimemload_24 & ((\Mux23~2_combout  & ((\my_reg[30][8]~q ))) # (!\Mux23~2_combout  & (\my_reg[26][8]~q )))) # (!dcifimemload_24 & (((\Mux23~2_combout ))))

	.dataa(\my_reg[26][8]~q ),
	.datab(\my_reg[30][8]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux23~2_combout ),
	.cin(gnd),
	.combout(\Mux23~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~3 .lut_mask = 16'hCFA0;
defparam \Mux23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N11
dffeas \my_reg[24][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][8] .is_wysiwyg = "true";
defparam \my_reg[24][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N19
dffeas \my_reg[28][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][8] .is_wysiwyg = "true";
defparam \my_reg[28][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N9
dffeas \my_reg[20][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][8] .is_wysiwyg = "true";
defparam \my_reg[20][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N13
dffeas \my_reg[16][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][8] .is_wysiwyg = "true";
defparam \my_reg[16][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N12
cycloneive_lcell_comb \Mux23~4 (
// Equation(s):
// \Mux23~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[20][8]~q )) # (!dcifimemload_23 & ((\my_reg[16][8]~q )))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[20][8]~q ),
	.datac(\my_reg[16][8]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux23~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~4 .lut_mask = 16'hEE50;
defparam \Mux23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N18
cycloneive_lcell_comb \Mux23~5 (
// Equation(s):
// \Mux23~5_combout  = (dcifimemload_24 & ((\Mux23~4_combout  & ((\my_reg[28][8]~q ))) # (!\Mux23~4_combout  & (\my_reg[24][8]~q )))) # (!dcifimemload_24 & (((\Mux23~4_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[24][8]~q ),
	.datac(\my_reg[28][8]~q ),
	.datad(\Mux23~4_combout ),
	.cin(gnd),
	.combout(\Mux23~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~5 .lut_mask = 16'hF588;
defparam \Mux23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N20
cycloneive_lcell_comb \Mux23~6 (
// Equation(s):
// \Mux23~6_combout  = (dcifimemload_22 & ((dcifimemload_21) # ((\Mux23~3_combout )))) # (!dcifimemload_22 & (!dcifimemload_21 & ((\Mux23~5_combout ))))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\Mux23~3_combout ),
	.datad(\Mux23~5_combout ),
	.cin(gnd),
	.combout(\Mux23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~6 .lut_mask = 16'hB9A8;
defparam \Mux23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N30
cycloneive_lcell_comb \Mux23~9 (
// Equation(s):
// \Mux23~9_combout  = (dcifimemload_21 & ((\Mux23~6_combout  & (\Mux23~8_combout )) # (!\Mux23~6_combout  & ((\Mux23~1_combout ))))) # (!dcifimemload_21 & (((\Mux23~6_combout ))))

	.dataa(\Mux23~8_combout ),
	.datab(dcifimemload_21),
	.datac(\Mux23~1_combout ),
	.datad(\Mux23~6_combout ),
	.cin(gnd),
	.combout(\Mux23~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~9 .lut_mask = 16'hBBC0;
defparam \Mux23~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N31
dffeas \my_reg[7][8] (
	.clk(CLK),
	.d(wdat25),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][8] .is_wysiwyg = "true";
defparam \my_reg[7][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N21
dffeas \my_reg[6][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][8] .is_wysiwyg = "true";
defparam \my_reg[6][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N10
cycloneive_lcell_comb \my_reg[5][8]~feeder (
// Equation(s):
// \my_reg[5][8]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat25),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[5][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[5][8]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[5][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N11
dffeas \my_reg[5][8] (
	.clk(CLK),
	.d(\my_reg[5][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][8] .is_wysiwyg = "true";
defparam \my_reg[5][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N28
cycloneive_lcell_comb \Mux23~10 (
// Equation(s):
// \Mux23~10_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\my_reg[5][8]~q ))) # (!dcifimemload_21 & (\my_reg[4][8]~q ))))

	.dataa(\my_reg[4][8]~q ),
	.datab(\my_reg[5][8]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux23~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~10 .lut_mask = 16'hFC0A;
defparam \Mux23~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N20
cycloneive_lcell_comb \Mux23~11 (
// Equation(s):
// \Mux23~11_combout  = (dcifimemload_22 & ((\Mux23~10_combout  & (\my_reg[7][8]~q )) # (!\Mux23~10_combout  & ((\my_reg[6][8]~q ))))) # (!dcifimemload_22 & (((\Mux23~10_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[7][8]~q ),
	.datac(\my_reg[6][8]~q ),
	.datad(\Mux23~10_combout ),
	.cin(gnd),
	.combout(\Mux23~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~11 .lut_mask = 16'hDDA0;
defparam \Mux23~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N14
cycloneive_lcell_comb \my_reg[14][8]~feeder (
// Equation(s):
// \my_reg[14][8]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat25),
	.cin(gnd),
	.combout(\my_reg[14][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[14][8]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[14][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N15
dffeas \my_reg[14][8] (
	.clk(CLK),
	.d(\my_reg[14][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][8] .is_wysiwyg = "true";
defparam \my_reg[14][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N5
dffeas \my_reg[13][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][8] .is_wysiwyg = "true";
defparam \my_reg[13][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N4
cycloneive_lcell_comb \Mux23~17 (
// Equation(s):
// \Mux23~17_combout  = (dcifimemload_21 & (((\my_reg[13][8]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\my_reg[12][8]~q  & ((!dcifimemload_22))))

	.dataa(\my_reg[12][8]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[13][8]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux23~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~17 .lut_mask = 16'hCCE2;
defparam \Mux23~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N28
cycloneive_lcell_comb \Mux23~18 (
// Equation(s):
// \Mux23~18_combout  = (\Mux23~17_combout  & ((\my_reg[15][8]~q ) # ((!dcifimemload_22)))) # (!\Mux23~17_combout  & (((\my_reg[14][8]~q  & dcifimemload_22))))

	.dataa(\my_reg[15][8]~q ),
	.datab(\my_reg[14][8]~q ),
	.datac(\Mux23~17_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux23~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~18 .lut_mask = 16'hACF0;
defparam \Mux23~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N21
dffeas \my_reg[1][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][8] .is_wysiwyg = "true";
defparam \my_reg[1][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N15
dffeas \my_reg[3][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][8] .is_wysiwyg = "true";
defparam \my_reg[3][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N14
cycloneive_lcell_comb \Mux23~14 (
// Equation(s):
// \Mux23~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][8]~q ))) # (!dcifimemload_22 & (\my_reg[1][8]~q ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[1][8]~q ),
	.datac(\my_reg[3][8]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux23~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~14 .lut_mask = 16'hA088;
defparam \Mux23~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N8
cycloneive_lcell_comb \Mux23~15 (
// Equation(s):
// \Mux23~15_combout  = (\Mux23~14_combout ) # ((\my_reg[2][8]~q  & (dcifimemload_22 & !dcifimemload_21)))

	.dataa(\my_reg[2][8]~q ),
	.datab(dcifimemload_22),
	.datac(dcifimemload_21),
	.datad(\Mux23~14_combout ),
	.cin(gnd),
	.combout(\Mux23~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~15 .lut_mask = 16'hFF08;
defparam \Mux23~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N23
dffeas \my_reg[11][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][8] .is_wysiwyg = "true";
defparam \my_reg[11][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N13
dffeas \my_reg[8][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][8] .is_wysiwyg = "true";
defparam \my_reg[8][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N12
cycloneive_lcell_comb \Mux23~12 (
// Equation(s):
// \Mux23~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][8]~q )) # (!dcifimemload_22 & ((\my_reg[8][8]~q )))))

	.dataa(\my_reg[10][8]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[8][8]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux23~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~12 .lut_mask = 16'hEE30;
defparam \Mux23~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N22
cycloneive_lcell_comb \Mux23~13 (
// Equation(s):
// \Mux23~13_combout  = (dcifimemload_21 & ((\Mux23~12_combout  & ((\my_reg[11][8]~q ))) # (!\Mux23~12_combout  & (\my_reg[9][8]~q )))) # (!dcifimemload_21 & (((\Mux23~12_combout ))))

	.dataa(\my_reg[9][8]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[11][8]~q ),
	.datad(\Mux23~12_combout ),
	.cin(gnd),
	.combout(\Mux23~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~13 .lut_mask = 16'hF388;
defparam \Mux23~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N2
cycloneive_lcell_comb \Mux23~16 (
// Equation(s):
// \Mux23~16_combout  = (dcifimemload_24 & ((dcifimemload_23) # ((\Mux23~13_combout )))) # (!dcifimemload_24 & (!dcifimemload_23 & (\Mux23~15_combout )))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux23~15_combout ),
	.datad(\Mux23~13_combout ),
	.cin(gnd),
	.combout(\Mux23~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~16 .lut_mask = 16'hBA98;
defparam \Mux23~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N28
cycloneive_lcell_comb \Mux23~19 (
// Equation(s):
// \Mux23~19_combout  = (dcifimemload_23 & ((\Mux23~16_combout  & ((\Mux23~18_combout ))) # (!\Mux23~16_combout  & (\Mux23~11_combout )))) # (!dcifimemload_23 & (((\Mux23~16_combout ))))

	.dataa(dcifimemload_23),
	.datab(\Mux23~11_combout ),
	.datac(\Mux23~18_combout ),
	.datad(\Mux23~16_combout ),
	.cin(gnd),
	.combout(\Mux23~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~19 .lut_mask = 16'hF588;
defparam \Mux23~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N15
dffeas \my_reg[12][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][8] .is_wysiwyg = "true";
defparam \my_reg[12][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N14
cycloneive_lcell_comb \Mux55~7 (
// Equation(s):
// \Mux55~7_combout  = (dcifimemload_17 & (dcifimemload_16)) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[13][8]~q ))) # (!dcifimemload_16 & (\my_reg[12][8]~q ))))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\my_reg[12][8]~q ),
	.datad(\my_reg[13][8]~q ),
	.cin(gnd),
	.combout(\Mux55~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~7 .lut_mask = 16'hDC98;
defparam \Mux55~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N17
dffeas \my_reg[15][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][8] .is_wysiwyg = "true";
defparam \my_reg[15][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N16
cycloneive_lcell_comb \Mux55~8 (
// Equation(s):
// \Mux55~8_combout  = (dcifimemload_17 & ((\Mux55~7_combout  & (\my_reg[15][8]~q )) # (!\Mux55~7_combout  & ((\my_reg[14][8]~q ))))) # (!dcifimemload_17 & (\Mux55~7_combout ))

	.dataa(dcifimemload_17),
	.datab(\Mux55~7_combout ),
	.datac(\my_reg[15][8]~q ),
	.datad(\my_reg[14][8]~q ),
	.cin(gnd),
	.combout(\Mux55~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~8 .lut_mask = 16'hE6C4;
defparam \Mux55~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N20
cycloneive_lcell_comb \Mux55~4 (
// Equation(s):
// \Mux55~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\my_reg[3][8]~q )) # (!dcifimemload_17 & ((\my_reg[1][8]~q )))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[3][8]~q ),
	.datac(\my_reg[1][8]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux55~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~4 .lut_mask = 16'h88A0;
defparam \Mux55~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N7
dffeas \my_reg[2][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][8] .is_wysiwyg = "true";
defparam \my_reg[2][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N6
cycloneive_lcell_comb \Mux55~5 (
// Equation(s):
// \Mux55~5_combout  = (\Mux55~4_combout ) # ((dcifimemload_17 & (\my_reg[2][8]~q  & !dcifimemload_16)))

	.dataa(dcifimemload_17),
	.datab(\Mux55~4_combout ),
	.datac(\my_reg[2][8]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux55~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~5 .lut_mask = 16'hCCEC;
defparam \Mux55~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N13
dffeas \my_reg[4][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][8] .is_wysiwyg = "true";
defparam \my_reg[4][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N12
cycloneive_lcell_comb \Mux55~2 (
// Equation(s):
// \Mux55~2_combout  = (dcifimemload_16 & ((\my_reg[5][8]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\my_reg[4][8]~q  & !dcifimemload_17))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[5][8]~q ),
	.datac(\my_reg[4][8]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux55~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~2 .lut_mask = 16'hAAD8;
defparam \Mux55~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N26
cycloneive_lcell_comb \Mux55~3 (
// Equation(s):
// \Mux55~3_combout  = (dcifimemload_17 & ((\Mux55~2_combout  & ((\my_reg[7][8]~q ))) # (!\Mux55~2_combout  & (\my_reg[6][8]~q )))) # (!dcifimemload_17 & (((\Mux55~2_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[6][8]~q ),
	.datac(\my_reg[7][8]~q ),
	.datad(\Mux55~2_combout ),
	.cin(gnd),
	.combout(\Mux55~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~3 .lut_mask = 16'hF588;
defparam \Mux55~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N22
cycloneive_lcell_comb \Mux55~6 (
// Equation(s):
// \Mux55~6_combout  = (dcifimemload_18 & ((dcifimemload_19) # ((\Mux55~3_combout )))) # (!dcifimemload_18 & (!dcifimemload_19 & (\Mux55~5_combout )))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux55~5_combout ),
	.datad(\Mux55~3_combout ),
	.cin(gnd),
	.combout(\Mux55~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~6 .lut_mask = 16'hBA98;
defparam \Mux55~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N18
cycloneive_lcell_comb \my_reg[9][8]~feeder (
// Equation(s):
// \my_reg[9][8]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat25),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[9][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[9][8]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[9][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N19
dffeas \my_reg[9][8] (
	.clk(CLK),
	.d(\my_reg[9][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][8] .is_wysiwyg = "true";
defparam \my_reg[9][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N13
dffeas \my_reg[10][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][8] .is_wysiwyg = "true";
defparam \my_reg[10][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N12
cycloneive_lcell_comb \Mux55~0 (
// Equation(s):
// \Mux55~0_combout  = (dcifimemload_17 & (((\my_reg[10][8]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\my_reg[8][8]~q  & ((!dcifimemload_16))))

	.dataa(\my_reg[8][8]~q ),
	.datab(dcifimemload_17),
	.datac(\my_reg[10][8]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux55~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~0 .lut_mask = 16'hCCE2;
defparam \Mux55~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N0
cycloneive_lcell_comb \Mux55~1 (
// Equation(s):
// \Mux55~1_combout  = (dcifimemload_16 & ((\Mux55~0_combout  & (\my_reg[11][8]~q )) # (!\Mux55~0_combout  & ((\my_reg[9][8]~q ))))) # (!dcifimemload_16 & (((\Mux55~0_combout ))))

	.dataa(\my_reg[11][8]~q ),
	.datab(\my_reg[9][8]~q ),
	.datac(dcifimemload_16),
	.datad(\Mux55~0_combout ),
	.cin(gnd),
	.combout(\Mux55~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~1 .lut_mask = 16'hAFC0;
defparam \Mux55~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N24
cycloneive_lcell_comb \my_reg[27][8]~feeder (
// Equation(s):
// \my_reg[27][8]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat25),
	.cin(gnd),
	.combout(\my_reg[27][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[27][8]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[27][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N25
dffeas \my_reg[27][8] (
	.clk(CLK),
	.d(\my_reg[27][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][8] .is_wysiwyg = "true";
defparam \my_reg[27][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N31
dffeas \my_reg[23][8] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][8] .is_wysiwyg = "true";
defparam \my_reg[23][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N30
cycloneive_lcell_comb \Mux55~17 (
// Equation(s):
// \Mux55~17_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[23][8]~q ))) # (!dcifimemload_18 & (\my_reg[19][8]~q ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[19][8]~q ),
	.datac(\my_reg[23][8]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux55~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~17 .lut_mask = 16'hFA44;
defparam \Mux55~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N12
cycloneive_lcell_comb \Mux55~18 (
// Equation(s):
// \Mux55~18_combout  = (dcifimemload_19 & ((\Mux55~17_combout  & ((\my_reg[31][8]~q ))) # (!\Mux55~17_combout  & (\my_reg[27][8]~q )))) # (!dcifimemload_19 & (((\Mux55~17_combout ))))

	.dataa(\my_reg[27][8]~q ),
	.datab(\my_reg[31][8]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux55~17_combout ),
	.cin(gnd),
	.combout(\Mux55~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~18 .lut_mask = 16'hCFA0;
defparam \Mux55~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N10
cycloneive_lcell_comb \Mux55~14 (
// Equation(s):
// \Mux55~14_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & (\my_reg[24][8]~q )) # (!dcifimemload_19 & ((\my_reg[16][8]~q )))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\my_reg[24][8]~q ),
	.datad(\my_reg[16][8]~q ),
	.cin(gnd),
	.combout(\Mux55~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~14 .lut_mask = 16'hD9C8;
defparam \Mux55~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N8
cycloneive_lcell_comb \Mux55~15 (
// Equation(s):
// \Mux55~15_combout  = (dcifimemload_18 & ((\Mux55~14_combout  & (\my_reg[28][8]~q )) # (!\Mux55~14_combout  & ((\my_reg[20][8]~q ))))) # (!dcifimemload_18 & (((\Mux55~14_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[28][8]~q ),
	.datac(\my_reg[20][8]~q ),
	.datad(\Mux55~14_combout ),
	.cin(gnd),
	.combout(\Mux55~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~15 .lut_mask = 16'hDDA0;
defparam \Mux55~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N0
cycloneive_lcell_comb \my_reg[26][8]~feeder (
// Equation(s):
// \my_reg[26][8]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat25),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[26][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[26][8]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[26][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y43_N1
dffeas \my_reg[26][8] (
	.clk(CLK),
	.d(\my_reg[26][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][8] .is_wysiwyg = "true";
defparam \my_reg[26][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N20
cycloneive_lcell_comb \Mux55~12 (
// Equation(s):
// \Mux55~12_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[26][8]~q ))) # (!dcifimemload_19 & (\my_reg[18][8]~q ))))

	.dataa(\my_reg[18][8]~q ),
	.datab(\my_reg[26][8]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux55~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~12 .lut_mask = 16'hFC0A;
defparam \Mux55~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N6
cycloneive_lcell_comb \Mux55~13 (
// Equation(s):
// \Mux55~13_combout  = (dcifimemload_18 & ((\Mux55~12_combout  & ((\my_reg[30][8]~q ))) # (!\Mux55~12_combout  & (\my_reg[22][8]~q )))) # (!dcifimemload_18 & (((\Mux55~12_combout ))))

	.dataa(\my_reg[22][8]~q ),
	.datab(\my_reg[30][8]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux55~12_combout ),
	.cin(gnd),
	.combout(\Mux55~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~13 .lut_mask = 16'hCFA0;
defparam \Mux55~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N4
cycloneive_lcell_comb \Mux55~16 (
// Equation(s):
// \Mux55~16_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux55~13_combout ))) # (!dcifimemload_17 & (\Mux55~15_combout ))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux55~15_combout ),
	.datad(\Mux55~13_combout ),
	.cin(gnd),
	.combout(\Mux55~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~16 .lut_mask = 16'hDC98;
defparam \Mux55~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N18
cycloneive_lcell_comb \my_reg[17][8]~feeder (
// Equation(s):
// \my_reg[17][8]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat25),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[17][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[17][8]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[17][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N19
dffeas \my_reg[17][8] (
	.clk(CLK),
	.d(\my_reg[17][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][8] .is_wysiwyg = "true";
defparam \my_reg[17][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N24
cycloneive_lcell_comb \Mux55~10 (
// Equation(s):
// \Mux55~10_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\my_reg[21][8]~q )) # (!dcifimemload_18 & ((\my_reg[17][8]~q )))))

	.dataa(\my_reg[21][8]~q ),
	.datab(\my_reg[17][8]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux55~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~10 .lut_mask = 16'hFA0C;
defparam \Mux55~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N18
cycloneive_lcell_comb \Mux55~11 (
// Equation(s):
// \Mux55~11_combout  = (dcifimemload_19 & ((\Mux55~10_combout  & (\my_reg[29][8]~q )) # (!\Mux55~10_combout  & ((\my_reg[25][8]~q ))))) # (!dcifimemload_19 & (((\Mux55~10_combout ))))

	.dataa(\my_reg[29][8]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[25][8]~q ),
	.datad(\Mux55~10_combout ),
	.cin(gnd),
	.combout(\Mux55~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~11 .lut_mask = 16'hBBC0;
defparam \Mux55~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N7
dffeas \my_reg[27][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][7] .is_wysiwyg = "true";
defparam \my_reg[27][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N11
dffeas \my_reg[31][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][7] .is_wysiwyg = "true";
defparam \my_reg[31][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N17
dffeas \my_reg[23][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][7] .is_wysiwyg = "true";
defparam \my_reg[23][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N16
cycloneive_lcell_comb \Mux24~7 (
// Equation(s):
// \Mux24~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\my_reg[23][7]~q ))) # (!dcifimemload_23 & (\my_reg[19][7]~q ))))

	.dataa(\my_reg[19][7]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[23][7]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux24~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~7 .lut_mask = 16'hFC22;
defparam \Mux24~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N10
cycloneive_lcell_comb \Mux24~8 (
// Equation(s):
// \Mux24~8_combout  = (dcifimemload_24 & ((\Mux24~7_combout  & ((\my_reg[31][7]~q ))) # (!\Mux24~7_combout  & (\my_reg[27][7]~q )))) # (!dcifimemload_24 & (((\Mux24~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[27][7]~q ),
	.datac(\my_reg[31][7]~q ),
	.datad(\Mux24~7_combout ),
	.cin(gnd),
	.combout(\Mux24~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~8 .lut_mask = 16'hF588;
defparam \Mux24~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N6
cycloneive_lcell_comb \my_reg[25][7]~feeder (
// Equation(s):
// \my_reg[25][7]~feeder_combout  = \wdat~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat26),
	.cin(gnd),
	.combout(\my_reg[25][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][7]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[25][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N7
dffeas \my_reg[25][7] (
	.clk(CLK),
	.d(\my_reg[25][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][7] .is_wysiwyg = "true";
defparam \my_reg[25][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N11
dffeas \my_reg[29][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][7] .is_wysiwyg = "true";
defparam \my_reg[29][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N20
cycloneive_lcell_comb \my_reg[17][7]~feeder (
// Equation(s):
// \my_reg[17][7]~feeder_combout  = \wdat~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat26),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[17][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[17][7]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[17][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N21
dffeas \my_reg[17][7] (
	.clk(CLK),
	.d(\my_reg[17][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][7] .is_wysiwyg = "true";
defparam \my_reg[17][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N1
dffeas \my_reg[21][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][7] .is_wysiwyg = "true";
defparam \my_reg[21][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N0
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\my_reg[21][7]~q ))) # (!dcifimemload_23 & (\my_reg[17][7]~q ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[17][7]~q ),
	.datac(\my_reg[21][7]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hFA44;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N12
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// \Mux24~1_combout  = (dcifimemload_24 & ((\Mux24~0_combout  & ((\my_reg[29][7]~q ))) # (!\Mux24~0_combout  & (\my_reg[25][7]~q )))) # (!dcifimemload_24 & (((\Mux24~0_combout ))))

	.dataa(\my_reg[25][7]~q ),
	.datab(\my_reg[29][7]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux24~0_combout ),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hCFA0;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N16
cycloneive_lcell_comb \my_reg[20][7]~feeder (
// Equation(s):
// \my_reg[20][7]~feeder_combout  = \wdat~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat26),
	.cin(gnd),
	.combout(\my_reg[20][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[20][7]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[20][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y31_N17
dffeas \my_reg[20][7] (
	.clk(CLK),
	.d(\my_reg[20][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][7] .is_wysiwyg = "true";
defparam \my_reg[20][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y42_N3
dffeas \my_reg[16][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][7] .is_wysiwyg = "true";
defparam \my_reg[16][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N4
cycloneive_lcell_comb \Mux24~4 (
// Equation(s):
// \Mux24~4_combout  = (dcifimemload_24 & ((\my_reg[24][7]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\my_reg[16][7]~q  & !dcifimemload_23))))

	.dataa(\my_reg[24][7]~q ),
	.datab(\my_reg[16][7]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~4 .lut_mask = 16'hF0AC;
defparam \Mux24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N6
cycloneive_lcell_comb \Mux24~5 (
// Equation(s):
// \Mux24~5_combout  = (\Mux24~4_combout  & ((\my_reg[28][7]~q ) # ((!dcifimemload_23)))) # (!\Mux24~4_combout  & (((\my_reg[20][7]~q  & dcifimemload_23))))

	.dataa(\my_reg[28][7]~q ),
	.datab(\my_reg[20][7]~q ),
	.datac(\Mux24~4_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~5 .lut_mask = 16'hACF0;
defparam \Mux24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N28
cycloneive_lcell_comb \my_reg[22][7]~feeder (
// Equation(s):
// \my_reg[22][7]~feeder_combout  = \wdat~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat26),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[22][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[22][7]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[22][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y43_N29
dffeas \my_reg[22][7] (
	.clk(CLK),
	.d(\my_reg[22][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][7] .is_wysiwyg = "true";
defparam \my_reg[22][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N14
cycloneive_lcell_comb \my_reg[26][7]~feeder (
// Equation(s):
// \my_reg[26][7]~feeder_combout  = \wdat~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat26),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[26][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[26][7]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[26][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y43_N15
dffeas \my_reg[26][7] (
	.clk(CLK),
	.d(\my_reg[26][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][7] .is_wysiwyg = "true";
defparam \my_reg[26][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N4
cycloneive_lcell_comb \Mux24~2 (
// Equation(s):
// \Mux24~2_combout  = (dcifimemload_24 & (((\my_reg[26][7]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\my_reg[18][7]~q  & ((!dcifimemload_23))))

	.dataa(\my_reg[18][7]~q ),
	.datab(\my_reg[26][7]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux24~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~2 .lut_mask = 16'hF0CA;
defparam \Mux24~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N18
cycloneive_lcell_comb \Mux24~3 (
// Equation(s):
// \Mux24~3_combout  = (\Mux24~2_combout  & ((\my_reg[30][7]~q ) # ((!dcifimemload_23)))) # (!\Mux24~2_combout  & (((\my_reg[22][7]~q  & dcifimemload_23))))

	.dataa(\my_reg[30][7]~q ),
	.datab(\my_reg[22][7]~q ),
	.datac(\Mux24~2_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux24~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~3 .lut_mask = 16'hACF0;
defparam \Mux24~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N0
cycloneive_lcell_comb \Mux24~6 (
// Equation(s):
// \Mux24~6_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux24~3_combout ))) # (!dcifimemload_22 & (\Mux24~5_combout ))))

	.dataa(\Mux24~5_combout ),
	.datab(dcifimemload_21),
	.datac(dcifimemload_22),
	.datad(\Mux24~3_combout ),
	.cin(gnd),
	.combout(\Mux24~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~6 .lut_mask = 16'hF2C2;
defparam \Mux24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N6
cycloneive_lcell_comb \my_reg[9][7]~feeder (
// Equation(s):
// \my_reg[9][7]~feeder_combout  = \wdat~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat26),
	.cin(gnd),
	.combout(\my_reg[9][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[9][7]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[9][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N7
dffeas \my_reg[9][7] (
	.clk(CLK),
	.d(\my_reg[9][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][7] .is_wysiwyg = "true";
defparam \my_reg[9][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N15
dffeas \my_reg[11][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][7] .is_wysiwyg = "true";
defparam \my_reg[11][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N1
dffeas \my_reg[8][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][7] .is_wysiwyg = "true";
defparam \my_reg[8][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N15
dffeas \my_reg[10][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][7] .is_wysiwyg = "true";
defparam \my_reg[10][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N14
cycloneive_lcell_comb \Mux24~10 (
// Equation(s):
// \Mux24~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[10][7]~q ))) # (!dcifimemload_22 & (\my_reg[8][7]~q ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[8][7]~q ),
	.datac(\my_reg[10][7]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux24~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~10 .lut_mask = 16'hFA44;
defparam \Mux24~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N12
cycloneive_lcell_comb \Mux24~11 (
// Equation(s):
// \Mux24~11_combout  = (dcifimemload_21 & ((\Mux24~10_combout  & ((\my_reg[11][7]~q ))) # (!\Mux24~10_combout  & (\my_reg[9][7]~q )))) # (!dcifimemload_21 & (((\Mux24~10_combout ))))

	.dataa(\my_reg[9][7]~q ),
	.datab(\my_reg[11][7]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux24~10_combout ),
	.cin(gnd),
	.combout(\Mux24~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~11 .lut_mask = 16'hCFA0;
defparam \Mux24~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N5
dffeas \my_reg[4][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][7] .is_wysiwyg = "true";
defparam \my_reg[4][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N4
cycloneive_lcell_comb \Mux24~12 (
// Equation(s):
// \Mux24~12_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\my_reg[5][7]~q )) # (!dcifimemload_21 & ((\my_reg[4][7]~q )))))

	.dataa(\my_reg[5][7]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[4][7]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux24~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~12 .lut_mask = 16'hEE30;
defparam \Mux24~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N27
dffeas \my_reg[7][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][7] .is_wysiwyg = "true";
defparam \my_reg[7][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N26
cycloneive_lcell_comb \Mux24~13 (
// Equation(s):
// \Mux24~13_combout  = (\Mux24~12_combout  & (((\my_reg[7][7]~q ) # (!dcifimemload_22)))) # (!\Mux24~12_combout  & (\my_reg[6][7]~q  & ((dcifimemload_22))))

	.dataa(\my_reg[6][7]~q ),
	.datab(\Mux24~12_combout ),
	.datac(\my_reg[7][7]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux24~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~13 .lut_mask = 16'hE2CC;
defparam \Mux24~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N25
dffeas \my_reg[2][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][7] .is_wysiwyg = "true";
defparam \my_reg[2][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N9
dffeas \my_reg[3][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][7] .is_wysiwyg = "true";
defparam \my_reg[3][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N8
cycloneive_lcell_comb \Mux24~14 (
// Equation(s):
// \Mux24~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][7]~q ))) # (!dcifimemload_22 & (\my_reg[1][7]~q ))))

	.dataa(\my_reg[1][7]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[3][7]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux24~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~14 .lut_mask = 16'hC088;
defparam \Mux24~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N20
cycloneive_lcell_comb \Mux24~15 (
// Equation(s):
// \Mux24~15_combout  = (\Mux24~14_combout ) # ((dcifimemload_22 & (\my_reg[2][7]~q  & !dcifimemload_21)))

	.dataa(dcifimemload_22),
	.datab(\my_reg[2][7]~q ),
	.datac(\Mux24~14_combout ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux24~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~15 .lut_mask = 16'hF0F8;
defparam \Mux24~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N26
cycloneive_lcell_comb \Mux24~16 (
// Equation(s):
// \Mux24~16_combout  = (dcifimemload_23 & ((dcifimemload_24) # ((\Mux24~13_combout )))) # (!dcifimemload_23 & (!dcifimemload_24 & ((\Mux24~15_combout ))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux24~13_combout ),
	.datad(\Mux24~15_combout ),
	.cin(gnd),
	.combout(\Mux24~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~16 .lut_mask = 16'hB9A8;
defparam \Mux24~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N27
dffeas \my_reg[13][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][7] .is_wysiwyg = "true";
defparam \my_reg[13][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N26
cycloneive_lcell_comb \Mux24~17 (
// Equation(s):
// \Mux24~17_combout  = (dcifimemload_21 & (((\my_reg[13][7]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\my_reg[12][7]~q  & ((!dcifimemload_22))))

	.dataa(\my_reg[12][7]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[13][7]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux24~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~17 .lut_mask = 16'hCCE2;
defparam \Mux24~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N26
cycloneive_lcell_comb \my_reg[15][7]~feeder (
// Equation(s):
// \my_reg[15][7]~feeder_combout  = \wdat~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat26),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[15][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[15][7]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[15][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N27
dffeas \my_reg[15][7] (
	.clk(CLK),
	.d(\my_reg[15][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][7] .is_wysiwyg = "true";
defparam \my_reg[15][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N31
dffeas \my_reg[14][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][7] .is_wysiwyg = "true";
defparam \my_reg[14][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N30
cycloneive_lcell_comb \Mux24~18 (
// Equation(s):
// \Mux24~18_combout  = (\Mux24~17_combout  & ((\my_reg[15][7]~q ) # ((!dcifimemload_22)))) # (!\Mux24~17_combout  & (((\my_reg[14][7]~q  & dcifimemload_22))))

	.dataa(\Mux24~17_combout ),
	.datab(\my_reg[15][7]~q ),
	.datac(\my_reg[14][7]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux24~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~18 .lut_mask = 16'hD8AA;
defparam \Mux24~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N23
dffeas \my_reg[12][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][7] .is_wysiwyg = "true";
defparam \my_reg[12][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N22
cycloneive_lcell_comb \Mux56~7 (
// Equation(s):
// \Mux56~7_combout  = (dcifimemload_17 & (dcifimemload_16)) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[13][7]~q ))) # (!dcifimemload_16 & (\my_reg[12][7]~q ))))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\my_reg[12][7]~q ),
	.datad(\my_reg[13][7]~q ),
	.cin(gnd),
	.combout(\Mux56~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~7 .lut_mask = 16'hDC98;
defparam \Mux56~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N14
cycloneive_lcell_comb \Mux56~8 (
// Equation(s):
// \Mux56~8_combout  = (dcifimemload_17 & ((\Mux56~7_combout  & (\my_reg[15][7]~q )) # (!\Mux56~7_combout  & ((\my_reg[14][7]~q ))))) # (!dcifimemload_17 & (((\Mux56~7_combout ))))

	.dataa(\my_reg[15][7]~q ),
	.datab(\my_reg[14][7]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux56~7_combout ),
	.cin(gnd),
	.combout(\Mux56~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~8 .lut_mask = 16'hAFC0;
defparam \Mux56~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N0
cycloneive_lcell_comb \Mux56~2 (
// Equation(s):
// \Mux56~2_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\my_reg[10][7]~q )) # (!dcifimemload_17 & ((\my_reg[8][7]~q )))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[10][7]~q ),
	.datac(\my_reg[8][7]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux56~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~2 .lut_mask = 16'hEE50;
defparam \Mux56~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N14
cycloneive_lcell_comb \Mux56~3 (
// Equation(s):
// \Mux56~3_combout  = (dcifimemload_16 & ((\Mux56~2_combout  & ((\my_reg[11][7]~q ))) # (!\Mux56~2_combout  & (\my_reg[9][7]~q )))) # (!dcifimemload_16 & (((\Mux56~2_combout ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[9][7]~q ),
	.datac(\my_reg[11][7]~q ),
	.datad(\Mux56~2_combout ),
	.cin(gnd),
	.combout(\Mux56~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~3 .lut_mask = 16'hF588;
defparam \Mux56~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N7
dffeas \my_reg[1][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][7] .is_wysiwyg = "true";
defparam \my_reg[1][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N6
cycloneive_lcell_comb \Mux56~4 (
// Equation(s):
// \Mux56~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\my_reg[3][7]~q )) # (!dcifimemload_17 & ((\my_reg[1][7]~q )))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[3][7]~q ),
	.datac(\my_reg[1][7]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux56~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~4 .lut_mask = 16'hD800;
defparam \Mux56~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N24
cycloneive_lcell_comb \Mux56~5 (
// Equation(s):
// \Mux56~5_combout  = (\Mux56~4_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \my_reg[2][7]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\my_reg[2][7]~q ),
	.datad(\Mux56~4_combout ),
	.cin(gnd),
	.combout(\Mux56~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~5 .lut_mask = 16'hFF20;
defparam \Mux56~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N8
cycloneive_lcell_comb \Mux56~6 (
// Equation(s):
// \Mux56~6_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\Mux56~3_combout )))) # (!dcifimemload_19 & (!dcifimemload_18 & ((\Mux56~5_combout ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux56~3_combout ),
	.datad(\Mux56~5_combout ),
	.cin(gnd),
	.combout(\Mux56~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~6 .lut_mask = 16'hB9A8;
defparam \Mux56~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y32_N9
dffeas \my_reg[6][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][7] .is_wysiwyg = "true";
defparam \my_reg[6][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N8
cycloneive_lcell_comb \my_reg[5][7]~feeder (
// Equation(s):
// \my_reg[5][7]~feeder_combout  = \wdat~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat26),
	.cin(gnd),
	.combout(\my_reg[5][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[5][7]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[5][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N9
dffeas \my_reg[5][7] (
	.clk(CLK),
	.d(\my_reg[5][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][7] .is_wysiwyg = "true";
defparam \my_reg[5][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N22
cycloneive_lcell_comb \Mux56~0 (
// Equation(s):
// \Mux56~0_combout  = (dcifimemload_16 & (((\my_reg[5][7]~q ) # (dcifimemload_17)))) # (!dcifimemload_16 & (\my_reg[4][7]~q  & ((!dcifimemload_17))))

	.dataa(\my_reg[4][7]~q ),
	.datab(\my_reg[5][7]~q ),
	.datac(dcifimemload_16),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux56~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~0 .lut_mask = 16'hF0CA;
defparam \Mux56~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N8
cycloneive_lcell_comb \Mux56~1 (
// Equation(s):
// \Mux56~1_combout  = (dcifimemload_17 & ((\Mux56~0_combout  & (\my_reg[7][7]~q )) # (!\Mux56~0_combout  & ((\my_reg[6][7]~q ))))) # (!dcifimemload_17 & (((\Mux56~0_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[7][7]~q ),
	.datac(\my_reg[6][7]~q ),
	.datad(\Mux56~0_combout ),
	.cin(gnd),
	.combout(\Mux56~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~1 .lut_mask = 16'hDDA0;
defparam \Mux56~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N6
cycloneive_lcell_comb \Mux56~17 (
// Equation(s):
// \Mux56~17_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[27][7]~q ))) # (!dcifimemload_19 & (\my_reg[19][7]~q ))))

	.dataa(\my_reg[19][7]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[27][7]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux56~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~17 .lut_mask = 16'hFC22;
defparam \Mux56~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N10
cycloneive_lcell_comb \Mux56~18 (
// Equation(s):
// \Mux56~18_combout  = (dcifimemload_18 & ((\Mux56~17_combout  & (\my_reg[31][7]~q )) # (!\Mux56~17_combout  & ((\my_reg[23][7]~q ))))) # (!dcifimemload_18 & (((\Mux56~17_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[31][7]~q ),
	.datac(\Mux56~17_combout ),
	.datad(\my_reg[23][7]~q ),
	.cin(gnd),
	.combout(\Mux56~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~18 .lut_mask = 16'hDAD0;
defparam \Mux56~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N24
cycloneive_lcell_comb \Mux56~10 (
// Equation(s):
// \Mux56~10_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[25][7]~q ))) # (!dcifimemload_19 & (\my_reg[17][7]~q ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[17][7]~q ),
	.datac(dcifimemload_19),
	.datad(\my_reg[25][7]~q ),
	.cin(gnd),
	.combout(\Mux56~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~10 .lut_mask = 16'hF4A4;
defparam \Mux56~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N10
cycloneive_lcell_comb \Mux56~11 (
// Equation(s):
// \Mux56~11_combout  = (dcifimemload_18 & ((\Mux56~10_combout  & ((\my_reg[29][7]~q ))) # (!\Mux56~10_combout  & (\my_reg[21][7]~q )))) # (!dcifimemload_18 & (((\Mux56~10_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[21][7]~q ),
	.datac(\my_reg[29][7]~q ),
	.datad(\Mux56~10_combout ),
	.cin(gnd),
	.combout(\Mux56~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~11 .lut_mask = 16'hF588;
defparam \Mux56~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N1
dffeas \my_reg[18][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][7] .is_wysiwyg = "true";
defparam \my_reg[18][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N0
cycloneive_lcell_comb \Mux56~12 (
// Equation(s):
// \Mux56~12_combout  = (dcifimemload_18 & ((\my_reg[22][7]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\my_reg[18][7]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[22][7]~q ),
	.datac(\my_reg[18][7]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux56~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~12 .lut_mask = 16'hAAD8;
defparam \Mux56~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N7
dffeas \my_reg[30][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][7] .is_wysiwyg = "true";
defparam \my_reg[30][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N6
cycloneive_lcell_comb \Mux56~13 (
// Equation(s):
// \Mux56~13_combout  = (\Mux56~12_combout  & (((\my_reg[30][7]~q ) # (!dcifimemload_19)))) # (!\Mux56~12_combout  & (\my_reg[26][7]~q  & ((dcifimemload_19))))

	.dataa(\my_reg[26][7]~q ),
	.datab(\Mux56~12_combout ),
	.datac(\my_reg[30][7]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux56~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~13 .lut_mask = 16'hE2CC;
defparam \Mux56~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y42_N1
dffeas \my_reg[28][7] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][7] .is_wysiwyg = "true";
defparam \my_reg[28][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N2
cycloneive_lcell_comb \Mux56~14 (
// Equation(s):
// \Mux56~14_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\my_reg[20][7]~q )) # (!dcifimemload_18 & ((\my_reg[16][7]~q )))))

	.dataa(\my_reg[20][7]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[16][7]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux56~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~14 .lut_mask = 16'hEE30;
defparam \Mux56~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N0
cycloneive_lcell_comb \Mux56~15 (
// Equation(s):
// \Mux56~15_combout  = (dcifimemload_19 & ((\Mux56~14_combout  & ((\my_reg[28][7]~q ))) # (!\Mux56~14_combout  & (\my_reg[24][7]~q )))) # (!dcifimemload_19 & (((\Mux56~14_combout ))))

	.dataa(\my_reg[24][7]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[28][7]~q ),
	.datad(\Mux56~14_combout ),
	.cin(gnd),
	.combout(\Mux56~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~15 .lut_mask = 16'hF388;
defparam \Mux56~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N20
cycloneive_lcell_comb \Mux56~16 (
// Equation(s):
// \Mux56~16_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\Mux56~13_combout )) # (!dcifimemload_17 & ((\Mux56~15_combout )))))

	.dataa(\Mux56~13_combout ),
	.datab(dcifimemload_16),
	.datac(dcifimemload_17),
	.datad(\Mux56~15_combout ),
	.cin(gnd),
	.combout(\Mux56~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~16 .lut_mask = 16'hE3E0;
defparam \Mux56~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N4
cycloneive_lcell_comb \my_reg[21][6]~feeder (
// Equation(s):
// \my_reg[21][6]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat27),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[21][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][6]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[21][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N5
dffeas \my_reg[21][6] (
	.clk(CLK),
	.d(\my_reg[21][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][6] .is_wysiwyg = "true";
defparam \my_reg[21][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N1
dffeas \my_reg[25][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][6] .is_wysiwyg = "true";
defparam \my_reg[25][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N0
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (dcifimemload_24 & (((\my_reg[25][6]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\my_reg[17][6]~q  & ((!dcifimemload_23))))

	.dataa(\my_reg[17][6]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[25][6]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hCCE2;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N5
dffeas \my_reg[29][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][6] .is_wysiwyg = "true";
defparam \my_reg[29][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N26
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (dcifimemload_23 & ((\Mux25~0_combout  & ((\my_reg[29][6]~q ))) # (!\Mux25~0_combout  & (\my_reg[21][6]~q )))) # (!dcifimemload_23 & (((\Mux25~0_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[21][6]~q ),
	.datac(\Mux25~0_combout ),
	.datad(\my_reg[29][6]~q ),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hF858;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N24
cycloneive_lcell_comb \my_reg[26][6]~feeder (
// Equation(s):
// \my_reg[26][6]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat27),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[26][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[26][6]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[26][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y43_N25
dffeas \my_reg[26][6] (
	.clk(CLK),
	.d(\my_reg[26][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][6] .is_wysiwyg = "true";
defparam \my_reg[26][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N22
cycloneive_lcell_comb \my_reg[22][6]~feeder (
// Equation(s):
// \my_reg[22][6]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat27),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[22][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[22][6]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[22][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y43_N23
dffeas \my_reg[22][6] (
	.clk(CLK),
	.d(\my_reg[22][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][6] .is_wysiwyg = "true";
defparam \my_reg[22][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N16
cycloneive_lcell_comb \Mux25~2 (
// Equation(s):
// \Mux25~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\my_reg[22][6]~q ))) # (!dcifimemload_23 & (\my_reg[18][6]~q ))))

	.dataa(\my_reg[18][6]~q ),
	.datab(\my_reg[22][6]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~2 .lut_mask = 16'hFC0A;
defparam \Mux25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N30
cycloneive_lcell_comb \Mux25~3 (
// Equation(s):
// \Mux25~3_combout  = (dcifimemload_24 & ((\Mux25~2_combout  & (\my_reg[30][6]~q )) # (!\Mux25~2_combout  & ((\my_reg[26][6]~q ))))) # (!dcifimemload_24 & (((\Mux25~2_combout ))))

	.dataa(\my_reg[30][6]~q ),
	.datab(\my_reg[26][6]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux25~2_combout ),
	.cin(gnd),
	.combout(\Mux25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~3 .lut_mask = 16'hAFC0;
defparam \Mux25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N24
cycloneive_lcell_comb \my_reg[24][6]~feeder (
// Equation(s):
// \my_reg[24][6]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat27),
	.cin(gnd),
	.combout(\my_reg[24][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[24][6]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[24][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y31_N25
dffeas \my_reg[24][6] (
	.clk(CLK),
	.d(\my_reg[24][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][6] .is_wysiwyg = "true";
defparam \my_reg[24][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y31_N19
dffeas \my_reg[20][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][6] .is_wysiwyg = "true";
defparam \my_reg[20][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N18
cycloneive_lcell_comb \Mux25~4 (
// Equation(s):
// \Mux25~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\my_reg[20][6]~q ))) # (!dcifimemload_23 & (\my_reg[16][6]~q ))))

	.dataa(\my_reg[16][6]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[20][6]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~4 .lut_mask = 16'hFC22;
defparam \Mux25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N12
cycloneive_lcell_comb \Mux25~5 (
// Equation(s):
// \Mux25~5_combout  = (dcifimemload_24 & ((\Mux25~4_combout  & (\my_reg[28][6]~q )) # (!\Mux25~4_combout  & ((\my_reg[24][6]~q ))))) # (!dcifimemload_24 & (((\Mux25~4_combout ))))

	.dataa(\my_reg[28][6]~q ),
	.datab(\my_reg[24][6]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux25~4_combout ),
	.cin(gnd),
	.combout(\Mux25~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~5 .lut_mask = 16'hAFC0;
defparam \Mux25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N22
cycloneive_lcell_comb \Mux25~6 (
// Equation(s):
// \Mux25~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & (\Mux25~3_combout )) # (!dcifimemload_22 & ((\Mux25~5_combout )))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux25~3_combout ),
	.datad(\Mux25~5_combout ),
	.cin(gnd),
	.combout(\Mux25~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~6 .lut_mask = 16'hD9C8;
defparam \Mux25~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N12
cycloneive_lcell_comb \my_reg[31][6]~feeder (
// Equation(s):
// \my_reg[31][6]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat27),
	.cin(gnd),
	.combout(\my_reg[31][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[31][6]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[31][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N13
dffeas \my_reg[31][6] (
	.clk(CLK),
	.d(\my_reg[31][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][6] .is_wysiwyg = "true";
defparam \my_reg[31][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N28
cycloneive_lcell_comb \my_reg[23][6]~feeder (
// Equation(s):
// \my_reg[23][6]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat27),
	.cin(gnd),
	.combout(\my_reg[23][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[23][6]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[23][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N29
dffeas \my_reg[23][6] (
	.clk(CLK),
	.d(\my_reg[23][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][6] .is_wysiwyg = "true";
defparam \my_reg[23][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N18
cycloneive_lcell_comb \my_reg[27][6]~feeder (
// Equation(s):
// \my_reg[27][6]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat27),
	.cin(gnd),
	.combout(\my_reg[27][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[27][6]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[27][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N19
dffeas \my_reg[27][6] (
	.clk(CLK),
	.d(\my_reg[27][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][6] .is_wysiwyg = "true";
defparam \my_reg[27][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N0
cycloneive_lcell_comb \Mux25~7 (
// Equation(s):
// \Mux25~7_combout  = (dcifimemload_24 & (((\my_reg[27][6]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\my_reg[19][6]~q  & ((!dcifimemload_23))))

	.dataa(\my_reg[19][6]~q ),
	.datab(\my_reg[27][6]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux25~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~7 .lut_mask = 16'hF0CA;
defparam \Mux25~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N26
cycloneive_lcell_comb \Mux25~8 (
// Equation(s):
// \Mux25~8_combout  = (dcifimemload_23 & ((\Mux25~7_combout  & (\my_reg[31][6]~q )) # (!\Mux25~7_combout  & ((\my_reg[23][6]~q ))))) # (!dcifimemload_23 & (((\Mux25~7_combout ))))

	.dataa(\my_reg[31][6]~q ),
	.datab(\my_reg[23][6]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux25~7_combout ),
	.cin(gnd),
	.combout(\Mux25~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~8 .lut_mask = 16'hAFC0;
defparam \Mux25~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N12
cycloneive_lcell_comb \my_reg[14][6]~feeder (
// Equation(s):
// \my_reg[14][6]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat27),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[14][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[14][6]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[14][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N13
dffeas \my_reg[14][6] (
	.clk(CLK),
	.d(\my_reg[14][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][6] .is_wysiwyg = "true";
defparam \my_reg[14][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N11
dffeas \my_reg[15][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][6] .is_wysiwyg = "true";
defparam \my_reg[15][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N16
cycloneive_lcell_comb \my_reg[13][6]~feeder (
// Equation(s):
// \my_reg[13][6]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat27),
	.cin(gnd),
	.combout(\my_reg[13][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[13][6]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[13][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N17
dffeas \my_reg[13][6] (
	.clk(CLK),
	.d(\my_reg[13][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][6] .is_wysiwyg = "true";
defparam \my_reg[13][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N30
cycloneive_lcell_comb \Mux25~17 (
// Equation(s):
// \Mux25~17_combout  = (dcifimemload_21 & (((\my_reg[13][6]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\my_reg[12][6]~q  & ((!dcifimemload_22))))

	.dataa(\my_reg[12][6]~q ),
	.datab(\my_reg[13][6]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux25~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~17 .lut_mask = 16'hF0CA;
defparam \Mux25~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N10
cycloneive_lcell_comb \Mux25~18 (
// Equation(s):
// \Mux25~18_combout  = (\Mux25~17_combout  & (((\my_reg[15][6]~q ) # (!dcifimemload_22)))) # (!\Mux25~17_combout  & (\my_reg[14][6]~q  & ((dcifimemload_22))))

	.dataa(\my_reg[14][6]~q ),
	.datab(\my_reg[15][6]~q ),
	.datac(\Mux25~17_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux25~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~18 .lut_mask = 16'hCAF0;
defparam \Mux25~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N10
cycloneive_lcell_comb \my_reg[7][6]~feeder (
// Equation(s):
// \my_reg[7][6]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat27),
	.cin(gnd),
	.combout(\my_reg[7][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[7][6]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[7][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y42_N11
dffeas \my_reg[7][6] (
	.clk(CLK),
	.d(\my_reg[7][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][6] .is_wysiwyg = "true";
defparam \my_reg[7][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N17
dffeas \my_reg[6][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][6] .is_wysiwyg = "true";
defparam \my_reg[6][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N0
cycloneive_lcell_comb \my_reg[4][6]~feeder (
// Equation(s):
// \my_reg[4][6]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat27),
	.cin(gnd),
	.combout(\my_reg[4][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[4][6]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[4][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y42_N1
dffeas \my_reg[4][6] (
	.clk(CLK),
	.d(\my_reg[4][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][6] .is_wysiwyg = "true";
defparam \my_reg[4][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N7
dffeas \my_reg[5][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][6] .is_wysiwyg = "true";
defparam \my_reg[5][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N6
cycloneive_lcell_comb \Mux25~10 (
// Equation(s):
// \Mux25~10_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\my_reg[5][6]~q ))) # (!dcifimemload_21 & (\my_reg[4][6]~q ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[4][6]~q ),
	.datac(\my_reg[5][6]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux25~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~10 .lut_mask = 16'hFA44;
defparam \Mux25~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N16
cycloneive_lcell_comb \Mux25~11 (
// Equation(s):
// \Mux25~11_combout  = (dcifimemload_22 & ((\Mux25~10_combout  & (\my_reg[7][6]~q )) # (!\Mux25~10_combout  & ((\my_reg[6][6]~q ))))) # (!dcifimemload_22 & (((\Mux25~10_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[7][6]~q ),
	.datac(\my_reg[6][6]~q ),
	.datad(\Mux25~10_combout ),
	.cin(gnd),
	.combout(\Mux25~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~11 .lut_mask = 16'hDDA0;
defparam \Mux25~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N3
dffeas \my_reg[10][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][6] .is_wysiwyg = "true";
defparam \my_reg[10][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N9
dffeas \my_reg[8][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][6] .is_wysiwyg = "true";
defparam \my_reg[8][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N8
cycloneive_lcell_comb \Mux25~12 (
// Equation(s):
// \Mux25~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][6]~q )) # (!dcifimemload_22 & ((\my_reg[8][6]~q )))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[10][6]~q ),
	.datac(\my_reg[8][6]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux25~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~12 .lut_mask = 16'hEE50;
defparam \Mux25~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N31
dffeas \my_reg[11][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][6] .is_wysiwyg = "true";
defparam \my_reg[11][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N30
cycloneive_lcell_comb \Mux25~13 (
// Equation(s):
// \Mux25~13_combout  = (\Mux25~12_combout  & (((\my_reg[11][6]~q ) # (!dcifimemload_21)))) # (!\Mux25~12_combout  & (\my_reg[9][6]~q  & ((dcifimemload_21))))

	.dataa(\my_reg[9][6]~q ),
	.datab(\Mux25~12_combout ),
	.datac(\my_reg[11][6]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux25~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~13 .lut_mask = 16'hE2CC;
defparam \Mux25~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N7
dffeas \my_reg[3][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][6] .is_wysiwyg = "true";
defparam \my_reg[3][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N28
cycloneive_lcell_comb \Mux25~14 (
// Equation(s):
// \Mux25~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][6]~q ))) # (!dcifimemload_22 & (\my_reg[1][6]~q ))))

	.dataa(\my_reg[1][6]~q ),
	.datab(\my_reg[3][6]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux25~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~14 .lut_mask = 16'hCA00;
defparam \Mux25~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N20
cycloneive_lcell_comb \Mux25~15 (
// Equation(s):
// \Mux25~15_combout  = (\Mux25~14_combout ) # ((\my_reg[2][6]~q  & (dcifimemload_22 & !dcifimemload_21)))

	.dataa(\my_reg[2][6]~q ),
	.datab(dcifimemload_22),
	.datac(dcifimemload_21),
	.datad(\Mux25~14_combout ),
	.cin(gnd),
	.combout(\Mux25~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~15 .lut_mask = 16'hFF08;
defparam \Mux25~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N2
cycloneive_lcell_comb \Mux25~16 (
// Equation(s):
// \Mux25~16_combout  = (dcifimemload_24 & ((dcifimemload_23) # ((\Mux25~13_combout )))) # (!dcifimemload_24 & (!dcifimemload_23 & ((\Mux25~15_combout ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux25~13_combout ),
	.datad(\Mux25~15_combout ),
	.cin(gnd),
	.combout(\Mux25~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~16 .lut_mask = 16'hB9A8;
defparam \Mux25~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N9
dffeas \my_reg[9][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][6] .is_wysiwyg = "true";
defparam \my_reg[9][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N2
cycloneive_lcell_comb \Mux57~0 (
// Equation(s):
// \Mux57~0_combout  = (dcifimemload_17 & (((\my_reg[10][6]~q ) # (dcifimemload_16)))) # (!dcifimemload_17 & (\my_reg[8][6]~q  & ((!dcifimemload_16))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[8][6]~q ),
	.datac(\my_reg[10][6]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux57~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~0 .lut_mask = 16'hAAE4;
defparam \Mux57~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N8
cycloneive_lcell_comb \Mux57~1 (
// Equation(s):
// \Mux57~1_combout  = (dcifimemload_16 & ((\Mux57~0_combout  & (\my_reg[11][6]~q )) # (!\Mux57~0_combout  & ((\my_reg[9][6]~q ))))) # (!dcifimemload_16 & (((\Mux57~0_combout ))))

	.dataa(\my_reg[11][6]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[9][6]~q ),
	.datad(\Mux57~0_combout ),
	.cin(gnd),
	.combout(\Mux57~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~1 .lut_mask = 16'hBBC0;
defparam \Mux57~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N8
cycloneive_lcell_comb \Mux57~2 (
// Equation(s):
// \Mux57~2_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][6]~q ))) # (!dcifimemload_16 & (\my_reg[4][6]~q ))))

	.dataa(\my_reg[4][6]~q ),
	.datab(\my_reg[5][6]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux57~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~2 .lut_mask = 16'hFC0A;
defparam \Mux57~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N2
cycloneive_lcell_comb \Mux57~3 (
// Equation(s):
// \Mux57~3_combout  = (dcifimemload_17 & ((\Mux57~2_combout  & (\my_reg[7][6]~q )) # (!\Mux57~2_combout  & ((\my_reg[6][6]~q ))))) # (!dcifimemload_17 & (((\Mux57~2_combout ))))

	.dataa(\my_reg[7][6]~q ),
	.datab(dcifimemload_17),
	.datac(\Mux57~2_combout ),
	.datad(\my_reg[6][6]~q ),
	.cin(gnd),
	.combout(\Mux57~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~3 .lut_mask = 16'hBCB0;
defparam \Mux57~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N27
dffeas \my_reg[2][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][6] .is_wysiwyg = "true";
defparam \my_reg[2][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N6
cycloneive_lcell_comb \Mux57~4 (
// Equation(s):
// \Mux57~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & ((\my_reg[3][6]~q ))) # (!dcifimemload_17 & (\my_reg[1][6]~q ))))

	.dataa(\my_reg[1][6]~q ),
	.datab(dcifimemload_16),
	.datac(\my_reg[3][6]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux57~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~4 .lut_mask = 16'hC088;
defparam \Mux57~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N26
cycloneive_lcell_comb \Mux57~5 (
// Equation(s):
// \Mux57~5_combout  = (\Mux57~4_combout ) # ((dcifimemload_17 & (!dcifimemload_16 & \my_reg[2][6]~q )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\my_reg[2][6]~q ),
	.datad(\Mux57~4_combout ),
	.cin(gnd),
	.combout(\Mux57~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~5 .lut_mask = 16'hFF20;
defparam \Mux57~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N30
cycloneive_lcell_comb \Mux57~6 (
// Equation(s):
// \Mux57~6_combout  = (dcifimemload_18 & ((dcifimemload_19) # ((\Mux57~3_combout )))) # (!dcifimemload_18 & (!dcifimemload_19 & ((\Mux57~5_combout ))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux57~3_combout ),
	.datad(\Mux57~5_combout ),
	.cin(gnd),
	.combout(\Mux57~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~6 .lut_mask = 16'hB9A8;
defparam \Mux57~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N29
dffeas \my_reg[12][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][6] .is_wysiwyg = "true";
defparam \my_reg[12][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N28
cycloneive_lcell_comb \Mux57~7 (
// Equation(s):
// \Mux57~7_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\my_reg[13][6]~q )) # (!dcifimemload_16 & ((\my_reg[12][6]~q )))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[13][6]~q ),
	.datac(\my_reg[12][6]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux57~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~7 .lut_mask = 16'hEE50;
defparam \Mux57~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N10
cycloneive_lcell_comb \Mux57~8 (
// Equation(s):
// \Mux57~8_combout  = (dcifimemload_17 & ((\Mux57~7_combout  & ((\my_reg[15][6]~q ))) # (!\Mux57~7_combout  & (\my_reg[14][6]~q )))) # (!dcifimemload_17 & (((\Mux57~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[14][6]~q ),
	.datac(\my_reg[15][6]~q ),
	.datad(\Mux57~7_combout ),
	.cin(gnd),
	.combout(\Mux57~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~8 .lut_mask = 16'hF588;
defparam \Mux57~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N2
cycloneive_lcell_comb \Mux57~10 (
// Equation(s):
// \Mux57~10_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[21][6]~q ))) # (!dcifimemload_18 & (\my_reg[17][6]~q ))))

	.dataa(\my_reg[17][6]~q ),
	.datab(\my_reg[21][6]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux57~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~10 .lut_mask = 16'hFC0A;
defparam \Mux57~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N4
cycloneive_lcell_comb \Mux57~11 (
// Equation(s):
// \Mux57~11_combout  = (dcifimemload_19 & ((\Mux57~10_combout  & ((\my_reg[29][6]~q ))) # (!\Mux57~10_combout  & (\my_reg[25][6]~q )))) # (!dcifimemload_19 & (((\Mux57~10_combout ))))

	.dataa(\my_reg[25][6]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[29][6]~q ),
	.datad(\Mux57~10_combout ),
	.cin(gnd),
	.combout(\Mux57~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~11 .lut_mask = 16'hF388;
defparam \Mux57~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N5
dffeas \my_reg[18][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][6] .is_wysiwyg = "true";
defparam \my_reg[18][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N4
cycloneive_lcell_comb \Mux57~12 (
// Equation(s):
// \Mux57~12_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\my_reg[26][6]~q )) # (!dcifimemload_19 & ((\my_reg[18][6]~q )))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[26][6]~q ),
	.datac(\my_reg[18][6]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux57~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~12 .lut_mask = 16'hEE50;
defparam \Mux57~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N23
dffeas \my_reg[30][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][6] .is_wysiwyg = "true";
defparam \my_reg[30][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N22
cycloneive_lcell_comb \Mux57~13 (
// Equation(s):
// \Mux57~13_combout  = (\Mux57~12_combout  & (((\my_reg[30][6]~q ) # (!dcifimemload_18)))) # (!\Mux57~12_combout  & (\my_reg[22][6]~q  & ((dcifimemload_18))))

	.dataa(\my_reg[22][6]~q ),
	.datab(\Mux57~12_combout ),
	.datac(\my_reg[30][6]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux57~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~13 .lut_mask = 16'hE2CC;
defparam \Mux57~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N21
dffeas \my_reg[16][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][6] .is_wysiwyg = "true";
defparam \my_reg[16][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N20
cycloneive_lcell_comb \Mux57~14 (
// Equation(s):
// \Mux57~14_combout  = (dcifimemload_19 & ((\my_reg[24][6]~q ) # ((dcifimemload_18)))) # (!dcifimemload_19 & (((\my_reg[16][6]~q  & !dcifimemload_18))))

	.dataa(\my_reg[24][6]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[16][6]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux57~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~14 .lut_mask = 16'hCCB8;
defparam \Mux57~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N19
dffeas \my_reg[28][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][6] .is_wysiwyg = "true";
defparam \my_reg[28][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N18
cycloneive_lcell_comb \Mux57~15 (
// Equation(s):
// \Mux57~15_combout  = (\Mux57~14_combout  & (((\my_reg[28][6]~q ) # (!dcifimemload_18)))) # (!\Mux57~14_combout  & (\my_reg[20][6]~q  & ((dcifimemload_18))))

	.dataa(\my_reg[20][6]~q ),
	.datab(\Mux57~14_combout ),
	.datac(\my_reg[28][6]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux57~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~15 .lut_mask = 16'hE2CC;
defparam \Mux57~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N8
cycloneive_lcell_comb \Mux57~16 (
// Equation(s):
// \Mux57~16_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & (\Mux57~13_combout )) # (!dcifimemload_17 & ((\Mux57~15_combout )))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux57~13_combout ),
	.datad(\Mux57~15_combout ),
	.cin(gnd),
	.combout(\Mux57~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~16 .lut_mask = 16'hD9C8;
defparam \Mux57~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N29
dffeas \my_reg[19][6] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][6] .is_wysiwyg = "true";
defparam \my_reg[19][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N28
cycloneive_lcell_comb \Mux57~17 (
// Equation(s):
// \Mux57~17_combout  = (dcifimemload_18 & ((\my_reg[23][6]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\my_reg[19][6]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[23][6]~q ),
	.datac(\my_reg[19][6]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux57~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~17 .lut_mask = 16'hAAD8;
defparam \Mux57~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N10
cycloneive_lcell_comb \Mux57~18 (
// Equation(s):
// \Mux57~18_combout  = (dcifimemload_19 & ((\Mux57~17_combout  & ((\my_reg[31][6]~q ))) # (!\Mux57~17_combout  & (\my_reg[27][6]~q )))) # (!dcifimemload_19 & (((\Mux57~17_combout ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[27][6]~q ),
	.datac(\Mux57~17_combout ),
	.datad(\my_reg[31][6]~q ),
	.cin(gnd),
	.combout(\Mux57~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~18 .lut_mask = 16'hF858;
defparam \Mux57~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N31
dffeas \my_reg[11][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][5] .is_wysiwyg = "true";
defparam \my_reg[11][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N5
dffeas \my_reg[9][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][5] .is_wysiwyg = "true";
defparam \my_reg[9][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N13
dffeas \my_reg[8][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][5] .is_wysiwyg = "true";
defparam \my_reg[8][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N26
cycloneive_lcell_comb \my_reg[10][5]~feeder (
// Equation(s):
// \my_reg[10][5]~feeder_combout  = \wdat~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat28),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[10][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[10][5]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[10][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N27
dffeas \my_reg[10][5] (
	.clk(CLK),
	.d(\my_reg[10][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][5] .is_wysiwyg = "true";
defparam \my_reg[10][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N16
cycloneive_lcell_comb \Mux26~10 (
// Equation(s):
// \Mux26~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[10][5]~q ))) # (!dcifimemload_22 & (\my_reg[8][5]~q ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[8][5]~q ),
	.datac(\my_reg[10][5]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux26~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~10 .lut_mask = 16'hFA44;
defparam \Mux26~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N4
cycloneive_lcell_comb \Mux26~11 (
// Equation(s):
// \Mux26~11_combout  = (dcifimemload_21 & ((\Mux26~10_combout  & (\my_reg[11][5]~q )) # (!\Mux26~10_combout  & ((\my_reg[9][5]~q ))))) # (!dcifimemload_21 & (((\Mux26~10_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[11][5]~q ),
	.datac(\my_reg[9][5]~q ),
	.datad(\Mux26~10_combout ),
	.cin(gnd),
	.combout(\Mux26~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~11 .lut_mask = 16'hDDA0;
defparam \Mux26~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N15
dffeas \my_reg[2][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][5] .is_wysiwyg = "true";
defparam \my_reg[2][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N25
dffeas \my_reg[1][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][5] .is_wysiwyg = "true";
defparam \my_reg[1][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N13
dffeas \my_reg[3][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][5] .is_wysiwyg = "true";
defparam \my_reg[3][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N12
cycloneive_lcell_comb \Mux26~14 (
// Equation(s):
// \Mux26~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][5]~q ))) # (!dcifimemload_22 & (\my_reg[1][5]~q ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[1][5]~q ),
	.datac(\my_reg[3][5]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux26~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~14 .lut_mask = 16'hA088;
defparam \Mux26~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N4
cycloneive_lcell_comb \Mux26~15 (
// Equation(s):
// \Mux26~15_combout  = (\Mux26~14_combout ) # ((!dcifimemload_21 & (\my_reg[2][5]~q  & dcifimemload_22)))

	.dataa(dcifimemload_21),
	.datab(\my_reg[2][5]~q ),
	.datac(dcifimemload_22),
	.datad(\Mux26~14_combout ),
	.cin(gnd),
	.combout(\Mux26~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~15 .lut_mask = 16'hFF40;
defparam \Mux26~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N11
dffeas \my_reg[7][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][5] .is_wysiwyg = "true";
defparam \my_reg[7][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N1
dffeas \my_reg[4][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][5] .is_wysiwyg = "true";
defparam \my_reg[4][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N0
cycloneive_lcell_comb \Mux26~12 (
// Equation(s):
// \Mux26~12_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\my_reg[5][5]~q )) # (!dcifimemload_21 & ((\my_reg[4][5]~q )))))

	.dataa(\my_reg[5][5]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[4][5]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux26~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~12 .lut_mask = 16'hEE30;
defparam \Mux26~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N10
cycloneive_lcell_comb \Mux26~13 (
// Equation(s):
// \Mux26~13_combout  = (dcifimemload_22 & ((\Mux26~12_combout  & ((\my_reg[7][5]~q ))) # (!\Mux26~12_combout  & (\my_reg[6][5]~q )))) # (!dcifimemload_22 & (((\Mux26~12_combout ))))

	.dataa(\my_reg[6][5]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[7][5]~q ),
	.datad(\Mux26~12_combout ),
	.cin(gnd),
	.combout(\Mux26~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~13 .lut_mask = 16'hF388;
defparam \Mux26~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N22
cycloneive_lcell_comb \Mux26~16 (
// Equation(s):
// \Mux26~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & ((\Mux26~13_combout ))) # (!dcifimemload_23 & (\Mux26~15_combout ))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux26~15_combout ),
	.datad(\Mux26~13_combout ),
	.cin(gnd),
	.combout(\Mux26~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~16 .lut_mask = 16'hDC98;
defparam \Mux26~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N20
cycloneive_lcell_comb \my_reg[14][5]~feeder (
// Equation(s):
// \my_reg[14][5]~feeder_combout  = \wdat~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat28),
	.cin(gnd),
	.combout(\my_reg[14][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[14][5]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[14][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N21
dffeas \my_reg[14][5] (
	.clk(CLK),
	.d(\my_reg[14][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][5] .is_wysiwyg = "true";
defparam \my_reg[14][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N9
dffeas \my_reg[13][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][5] .is_wysiwyg = "true";
defparam \my_reg[13][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N8
cycloneive_lcell_comb \Mux26~17 (
// Equation(s):
// \Mux26~17_combout  = (dcifimemload_21 & (((\my_reg[13][5]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\my_reg[12][5]~q  & ((!dcifimemload_22))))

	.dataa(\my_reg[12][5]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[13][5]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux26~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~17 .lut_mask = 16'hCCE2;
defparam \Mux26~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N6
cycloneive_lcell_comb \Mux26~18 (
// Equation(s):
// \Mux26~18_combout  = (dcifimemload_22 & ((\Mux26~17_combout  & (\my_reg[15][5]~q )) # (!\Mux26~17_combout  & ((\my_reg[14][5]~q ))))) # (!dcifimemload_22 & (((\Mux26~17_combout ))))

	.dataa(\my_reg[15][5]~q ),
	.datab(\my_reg[14][5]~q ),
	.datac(dcifimemload_22),
	.datad(\Mux26~17_combout ),
	.cin(gnd),
	.combout(\Mux26~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~18 .lut_mask = 16'hAFC0;
defparam \Mux26~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N12
cycloneive_lcell_comb \Mux26~19 (
// Equation(s):
// \Mux26~19_combout  = (dcifimemload_24 & ((\Mux26~16_combout  & ((\Mux26~18_combout ))) # (!\Mux26~16_combout  & (\Mux26~11_combout )))) # (!dcifimemload_24 & (((\Mux26~16_combout ))))

	.dataa(\Mux26~11_combout ),
	.datab(dcifimemload_24),
	.datac(\Mux26~16_combout ),
	.datad(\Mux26~18_combout ),
	.cin(gnd),
	.combout(\Mux26~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~19 .lut_mask = 16'hF838;
defparam \Mux26~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y34_N1
dffeas \my_reg[27][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][5] .is_wysiwyg = "true";
defparam \my_reg[27][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N7
dffeas \my_reg[19][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][5] .is_wysiwyg = "true";
defparam \my_reg[19][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N6
cycloneive_lcell_comb \Mux26~7 (
// Equation(s):
// \Mux26~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[23][5]~q )) # (!dcifimemload_23 & ((\my_reg[19][5]~q )))))

	.dataa(\my_reg[23][5]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[19][5]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux26~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~7 .lut_mask = 16'hEE30;
defparam \Mux26~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N0
cycloneive_lcell_comb \Mux26~8 (
// Equation(s):
// \Mux26~8_combout  = (dcifimemload_24 & ((\Mux26~7_combout  & (\my_reg[31][5]~q )) # (!\Mux26~7_combout  & ((\my_reg[27][5]~q ))))) # (!dcifimemload_24 & (((\Mux26~7_combout ))))

	.dataa(\my_reg[31][5]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[27][5]~q ),
	.datad(\Mux26~7_combout ),
	.cin(gnd),
	.combout(\Mux26~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~8 .lut_mask = 16'hBBC0;
defparam \Mux26~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N31
dffeas \my_reg[29][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][5] .is_wysiwyg = "true";
defparam \my_reg[29][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N10
cycloneive_lcell_comb \my_reg[21][5]~feeder (
// Equation(s):
// \my_reg[21][5]~feeder_combout  = \wdat~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat28),
	.cin(gnd),
	.combout(\my_reg[21][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][5]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[21][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y31_N11
dffeas \my_reg[21][5] (
	.clk(CLK),
	.d(\my_reg[21][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][5] .is_wysiwyg = "true";
defparam \my_reg[21][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N24
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (dcifimemload_23 & (((\my_reg[21][5]~q ) # (dcifimemload_24)))) # (!dcifimemload_23 & (\my_reg[17][5]~q  & ((!dcifimemload_24))))

	.dataa(\my_reg[17][5]~q ),
	.datab(\my_reg[21][5]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hF0CA;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N30
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (dcifimemload_24 & ((\Mux26~0_combout  & ((\my_reg[29][5]~q ))) # (!\Mux26~0_combout  & (\my_reg[25][5]~q )))) # (!dcifimemload_24 & (((\Mux26~0_combout ))))

	.dataa(\my_reg[25][5]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[29][5]~q ),
	.datad(\Mux26~0_combout ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hF388;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N26
cycloneive_lcell_comb \my_reg[28][5]~feeder (
// Equation(s):
// \my_reg[28][5]~feeder_combout  = \wdat~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat28),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[28][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[28][5]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[28][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y32_N27
dffeas \my_reg[28][5] (
	.clk(CLK),
	.d(\my_reg[28][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][5] .is_wysiwyg = "true";
defparam \my_reg[28][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y31_N15
dffeas \my_reg[20][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][5] .is_wysiwyg = "true";
defparam \my_reg[20][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N0
cycloneive_lcell_comb \my_reg[16][5]~feeder (
// Equation(s):
// \my_reg[16][5]~feeder_combout  = \wdat~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat28),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[16][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[16][5]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[16][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y32_N1
dffeas \my_reg[16][5] (
	.clk(CLK),
	.d(\my_reg[16][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][5] .is_wysiwyg = "true";
defparam \my_reg[16][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N10
cycloneive_lcell_comb \Mux26~4 (
// Equation(s):
// \Mux26~4_combout  = (dcifimemload_24 & ((\my_reg[24][5]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\my_reg[16][5]~q  & !dcifimemload_23))))

	.dataa(\my_reg[24][5]~q ),
	.datab(\my_reg[16][5]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~4 .lut_mask = 16'hF0AC;
defparam \Mux26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N14
cycloneive_lcell_comb \Mux26~5 (
// Equation(s):
// \Mux26~5_combout  = (dcifimemload_23 & ((\Mux26~4_combout  & (\my_reg[28][5]~q )) # (!\Mux26~4_combout  & ((\my_reg[20][5]~q ))))) # (!dcifimemload_23 & (((\Mux26~4_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[28][5]~q ),
	.datac(\my_reg[20][5]~q ),
	.datad(\Mux26~4_combout ),
	.cin(gnd),
	.combout(\Mux26~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~5 .lut_mask = 16'hDDA0;
defparam \Mux26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N15
dffeas \my_reg[30][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][5] .is_wysiwyg = "true";
defparam \my_reg[30][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N29
dffeas \my_reg[18][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][5] .is_wysiwyg = "true";
defparam \my_reg[18][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N8
cycloneive_lcell_comb \Mux26~2 (
// Equation(s):
// \Mux26~2_combout  = (dcifimemload_24 & ((\my_reg[26][5]~q ) # ((dcifimemload_23)))) # (!dcifimemload_24 & (((\my_reg[18][5]~q  & !dcifimemload_23))))

	.dataa(\my_reg[26][5]~q ),
	.datab(\my_reg[18][5]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~2 .lut_mask = 16'hF0AC;
defparam \Mux26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N22
cycloneive_lcell_comb \Mux26~3 (
// Equation(s):
// \Mux26~3_combout  = (\Mux26~2_combout  & (((\my_reg[30][5]~q ) # (!dcifimemload_23)))) # (!\Mux26~2_combout  & (\my_reg[22][5]~q  & ((dcifimemload_23))))

	.dataa(\my_reg[22][5]~q ),
	.datab(\my_reg[30][5]~q ),
	.datac(\Mux26~2_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~3 .lut_mask = 16'hCAF0;
defparam \Mux26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N28
cycloneive_lcell_comb \Mux26~6 (
// Equation(s):
// \Mux26~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux26~3_combout ))) # (!dcifimemload_22 & (\Mux26~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux26~5_combout ),
	.datad(\Mux26~3_combout ),
	.cin(gnd),
	.combout(\Mux26~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~6 .lut_mask = 16'hDC98;
defparam \Mux26~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N2
cycloneive_lcell_comb \Mux26~9 (
// Equation(s):
// \Mux26~9_combout  = (dcifimemload_21 & ((\Mux26~6_combout  & (\Mux26~8_combout )) # (!\Mux26~6_combout  & ((\Mux26~1_combout ))))) # (!dcifimemload_21 & (((\Mux26~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux26~8_combout ),
	.datac(\Mux26~1_combout ),
	.datad(\Mux26~6_combout ),
	.cin(gnd),
	.combout(\Mux26~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~9 .lut_mask = 16'hDDA0;
defparam \Mux26~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y32_N9
dffeas \my_reg[6][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][5] .is_wysiwyg = "true";
defparam \my_reg[6][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y32_N3
dffeas \my_reg[5][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][5] .is_wysiwyg = "true";
defparam \my_reg[5][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N2
cycloneive_lcell_comb \Mux58~0 (
// Equation(s):
// \Mux58~0_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][5]~q ))) # (!dcifimemload_16 & (\my_reg[4][5]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[4][5]~q ),
	.datac(\my_reg[5][5]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux58~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~0 .lut_mask = 16'hFA44;
defparam \Mux58~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N8
cycloneive_lcell_comb \Mux58~1 (
// Equation(s):
// \Mux58~1_combout  = (dcifimemload_17 & ((\Mux58~0_combout  & (\my_reg[7][5]~q )) # (!\Mux58~0_combout  & ((\my_reg[6][5]~q ))))) # (!dcifimemload_17 & (((\Mux58~0_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[7][5]~q ),
	.datac(\my_reg[6][5]~q ),
	.datad(\Mux58~0_combout ),
	.cin(gnd),
	.combout(\Mux58~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~1 .lut_mask = 16'hDDA0;
defparam \Mux58~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N31
dffeas \my_reg[15][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][5] .is_wysiwyg = "true";
defparam \my_reg[15][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N1
dffeas \my_reg[12][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][5] .is_wysiwyg = "true";
defparam \my_reg[12][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N0
cycloneive_lcell_comb \Mux58~7 (
// Equation(s):
// \Mux58~7_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\my_reg[13][5]~q )) # (!dcifimemload_16 & ((\my_reg[12][5]~q )))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[13][5]~q ),
	.datac(\my_reg[12][5]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux58~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~7 .lut_mask = 16'hEE50;
defparam \Mux58~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N30
cycloneive_lcell_comb \Mux58~8 (
// Equation(s):
// \Mux58~8_combout  = (dcifimemload_17 & ((\Mux58~7_combout  & ((\my_reg[15][5]~q ))) # (!\Mux58~7_combout  & (\my_reg[14][5]~q )))) # (!dcifimemload_17 & (((\Mux58~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[14][5]~q ),
	.datac(\my_reg[15][5]~q ),
	.datad(\Mux58~7_combout ),
	.cin(gnd),
	.combout(\Mux58~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~8 .lut_mask = 16'hF588;
defparam \Mux58~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N24
cycloneive_lcell_comb \Mux58~4 (
// Equation(s):
// \Mux58~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\my_reg[3][5]~q )) # (!dcifimemload_17 & ((\my_reg[1][5]~q )))))

	.dataa(\my_reg[3][5]~q ),
	.datab(dcifimemload_17),
	.datac(\my_reg[1][5]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux58~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~4 .lut_mask = 16'hB800;
defparam \Mux58~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N14
cycloneive_lcell_comb \Mux58~5 (
// Equation(s):
// \Mux58~5_combout  = (\Mux58~4_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \my_reg[2][5]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\my_reg[2][5]~q ),
	.datad(\Mux58~4_combout ),
	.cin(gnd),
	.combout(\Mux58~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~5 .lut_mask = 16'hFF40;
defparam \Mux58~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N12
cycloneive_lcell_comb \Mux58~2 (
// Equation(s):
// \Mux58~2_combout  = (dcifimemload_17 & ((\my_reg[10][5]~q ) # ((dcifimemload_16)))) # (!dcifimemload_17 & (((\my_reg[8][5]~q  & !dcifimemload_16))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[10][5]~q ),
	.datac(\my_reg[8][5]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux58~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~2 .lut_mask = 16'hAAD8;
defparam \Mux58~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N30
cycloneive_lcell_comb \Mux58~3 (
// Equation(s):
// \Mux58~3_combout  = (dcifimemload_16 & ((\Mux58~2_combout  & ((\my_reg[11][5]~q ))) # (!\Mux58~2_combout  & (\my_reg[9][5]~q )))) # (!dcifimemload_16 & (((\Mux58~2_combout ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[9][5]~q ),
	.datac(\my_reg[11][5]~q ),
	.datad(\Mux58~2_combout ),
	.cin(gnd),
	.combout(\Mux58~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~3 .lut_mask = 16'hF588;
defparam \Mux58~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N28
cycloneive_lcell_comb \Mux58~6 (
// Equation(s):
// \Mux58~6_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & ((\Mux58~3_combout ))) # (!dcifimemload_19 & (\Mux58~5_combout ))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux58~5_combout ),
	.datad(\Mux58~3_combout ),
	.cin(gnd),
	.combout(\Mux58~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~6 .lut_mask = 16'hDC98;
defparam \Mux58~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N12
cycloneive_lcell_comb \Mux58~17 (
// Equation(s):
// \Mux58~17_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\my_reg[27][5]~q )) # (!dcifimemload_19 & ((\my_reg[19][5]~q )))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[27][5]~q ),
	.datac(dcifimemload_19),
	.datad(\my_reg[19][5]~q ),
	.cin(gnd),
	.combout(\Mux58~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~17 .lut_mask = 16'hE5E0;
defparam \Mux58~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N4
cycloneive_lcell_comb \my_reg[23][5]~feeder (
// Equation(s):
// \my_reg[23][5]~feeder_combout  = \wdat~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat28),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[23][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[23][5]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[23][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N5
dffeas \my_reg[23][5] (
	.clk(CLK),
	.d(\my_reg[23][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][5] .is_wysiwyg = "true";
defparam \my_reg[23][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N19
dffeas \my_reg[31][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][5] .is_wysiwyg = "true";
defparam \my_reg[31][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N18
cycloneive_lcell_comb \Mux58~18 (
// Equation(s):
// \Mux58~18_combout  = (\Mux58~17_combout  & (((\my_reg[31][5]~q ) # (!dcifimemload_18)))) # (!\Mux58~17_combout  & (\my_reg[23][5]~q  & ((dcifimemload_18))))

	.dataa(\Mux58~17_combout ),
	.datab(\my_reg[23][5]~q ),
	.datac(\my_reg[31][5]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux58~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~18 .lut_mask = 16'hE4AA;
defparam \Mux58~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N0
cycloneive_lcell_comb \my_reg[24][5]~feeder (
// Equation(s):
// \my_reg[24][5]~feeder_combout  = \wdat~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat28),
	.cin(gnd),
	.combout(\my_reg[24][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[24][5]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[24][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y31_N1
dffeas \my_reg[24][5] (
	.clk(CLK),
	.d(\my_reg[24][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][5] .is_wysiwyg = "true";
defparam \my_reg[24][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N2
cycloneive_lcell_comb \Mux58~14 (
// Equation(s):
// \Mux58~14_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[20][5]~q ))) # (!dcifimemload_18 & (\my_reg[16][5]~q ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[16][5]~q ),
	.datac(dcifimemload_18),
	.datad(\my_reg[20][5]~q ),
	.cin(gnd),
	.combout(\Mux58~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~14 .lut_mask = 16'hF4A4;
defparam \Mux58~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N12
cycloneive_lcell_comb \Mux58~15 (
// Equation(s):
// \Mux58~15_combout  = (dcifimemload_19 & ((\Mux58~14_combout  & (\my_reg[28][5]~q )) # (!\Mux58~14_combout  & ((\my_reg[24][5]~q ))))) # (!dcifimemload_19 & (((\Mux58~14_combout ))))

	.dataa(\my_reg[28][5]~q ),
	.datab(\my_reg[24][5]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux58~14_combout ),
	.cin(gnd),
	.combout(\Mux58~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~15 .lut_mask = 16'hAFC0;
defparam \Mux58~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N12
cycloneive_lcell_comb \my_reg[22][5]~feeder (
// Equation(s):
// \my_reg[22][5]~feeder_combout  = \wdat~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat28),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[22][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[22][5]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[22][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y43_N13
dffeas \my_reg[22][5] (
	.clk(CLK),
	.d(\my_reg[22][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][5] .is_wysiwyg = "true";
defparam \my_reg[22][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N28
cycloneive_lcell_comb \Mux58~12 (
// Equation(s):
// \Mux58~12_combout  = (dcifimemload_18 & ((\my_reg[22][5]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\my_reg[18][5]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[22][5]~q ),
	.datac(\my_reg[18][5]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux58~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~12 .lut_mask = 16'hAAD8;
defparam \Mux58~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N14
cycloneive_lcell_comb \Mux58~13 (
// Equation(s):
// \Mux58~13_combout  = (\Mux58~12_combout  & (((\my_reg[30][5]~q ) # (!dcifimemload_19)))) # (!\Mux58~12_combout  & (\my_reg[26][5]~q  & ((dcifimemload_19))))

	.dataa(\my_reg[26][5]~q ),
	.datab(\Mux58~12_combout ),
	.datac(\my_reg[30][5]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux58~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~13 .lut_mask = 16'hE2CC;
defparam \Mux58~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N30
cycloneive_lcell_comb \Mux58~16 (
// Equation(s):
// \Mux58~16_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux58~13_combout ))) # (!dcifimemload_17 & (\Mux58~15_combout ))))

	.dataa(\Mux58~15_combout ),
	.datab(dcifimemload_16),
	.datac(dcifimemload_17),
	.datad(\Mux58~13_combout ),
	.cin(gnd),
	.combout(\Mux58~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~16 .lut_mask = 16'hF2C2;
defparam \Mux58~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N9
dffeas \my_reg[17][5] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][5] .is_wysiwyg = "true";
defparam \my_reg[17][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N8
cycloneive_lcell_comb \Mux58~10 (
// Equation(s):
// \Mux58~10_combout  = (dcifimemload_19 & ((\my_reg[25][5]~q ) # ((dcifimemload_18)))) # (!dcifimemload_19 & (((\my_reg[17][5]~q  & !dcifimemload_18))))

	.dataa(\my_reg[25][5]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[17][5]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux58~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~10 .lut_mask = 16'hCCB8;
defparam \Mux58~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N22
cycloneive_lcell_comb \Mux58~11 (
// Equation(s):
// \Mux58~11_combout  = (\Mux58~10_combout  & (((\my_reg[29][5]~q ) # (!dcifimemload_18)))) # (!\Mux58~10_combout  & (\my_reg[21][5]~q  & ((dcifimemload_18))))

	.dataa(\my_reg[21][5]~q ),
	.datab(\my_reg[29][5]~q ),
	.datac(\Mux58~10_combout ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux58~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~11 .lut_mask = 16'hCAF0;
defparam \Mux58~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N0
cycloneive_lcell_comb \my_reg[29][4]~feeder (
// Equation(s):
// \my_reg[29][4]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat29),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[29][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[29][4]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[29][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N1
dffeas \my_reg[29][4] (
	.clk(CLK),
	.d(\my_reg[29][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][4] .is_wysiwyg = "true";
defparam \my_reg[29][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N0
cycloneive_lcell_comb \my_reg[21][4]~feeder (
// Equation(s):
// \my_reg[21][4]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat29),
	.cin(gnd),
	.combout(\my_reg[21][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][4]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[21][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N1
dffeas \my_reg[21][4] (
	.clk(CLK),
	.d(\my_reg[21][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][4] .is_wysiwyg = "true";
defparam \my_reg[21][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N20
cycloneive_lcell_comb \my_reg[25][4]~feeder (
// Equation(s):
// \my_reg[25][4]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat29),
	.cin(gnd),
	.combout(\my_reg[25][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][4]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[25][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N21
dffeas \my_reg[25][4] (
	.clk(CLK),
	.d(\my_reg[25][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][4] .is_wysiwyg = "true";
defparam \my_reg[25][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N14
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & ((\my_reg[25][4]~q ))) # (!dcifimemload_24 & (\my_reg[17][4]~q ))))

	.dataa(\my_reg[17][4]~q ),
	.datab(\my_reg[25][4]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hFC0A;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N18
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// \Mux27~1_combout  = (dcifimemload_23 & ((\Mux27~0_combout  & (\my_reg[29][4]~q )) # (!\Mux27~0_combout  & ((\my_reg[21][4]~q ))))) # (!dcifimemload_23 & (((\Mux27~0_combout ))))

	.dataa(\my_reg[29][4]~q ),
	.datab(\my_reg[21][4]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux27~0_combout ),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hAFC0;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N22
cycloneive_lcell_comb \my_reg[31][4]~feeder (
// Equation(s):
// \my_reg[31][4]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat29),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[31][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[31][4]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[31][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N23
dffeas \my_reg[31][4] (
	.clk(CLK),
	.d(\my_reg[31][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][4] .is_wysiwyg = "true";
defparam \my_reg[31][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N26
cycloneive_lcell_comb \my_reg[23][4]~feeder (
// Equation(s):
// \my_reg[23][4]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat29),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[23][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[23][4]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[23][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N27
dffeas \my_reg[23][4] (
	.clk(CLK),
	.d(\my_reg[23][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][4] .is_wysiwyg = "true";
defparam \my_reg[23][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N20
cycloneive_lcell_comb \my_reg[19][4]~feeder (
// Equation(s):
// \my_reg[19][4]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat29),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[19][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[19][4]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[19][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N21
dffeas \my_reg[19][4] (
	.clk(CLK),
	.d(\my_reg[19][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][4] .is_wysiwyg = "true";
defparam \my_reg[19][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y36_N31
dffeas \my_reg[27][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][4] .is_wysiwyg = "true";
defparam \my_reg[27][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N30
cycloneive_lcell_comb \Mux27~7 (
// Equation(s):
// \Mux27~7_combout  = (dcifimemload_24 & (((\my_reg[27][4]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\my_reg[19][4]~q  & ((!dcifimemload_23))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[19][4]~q ),
	.datac(\my_reg[27][4]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux27~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~7 .lut_mask = 16'hAAE4;
defparam \Mux27~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N26
cycloneive_lcell_comb \Mux27~8 (
// Equation(s):
// \Mux27~8_combout  = (\Mux27~7_combout  & ((\my_reg[31][4]~q ) # ((!dcifimemload_23)))) # (!\Mux27~7_combout  & (((\my_reg[23][4]~q  & dcifimemload_23))))

	.dataa(\my_reg[31][4]~q ),
	.datab(\my_reg[23][4]~q ),
	.datac(\Mux27~7_combout ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux27~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~8 .lut_mask = 16'hACF0;
defparam \Mux27~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y31_N29
dffeas \my_reg[24][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][4] .is_wysiwyg = "true";
defparam \my_reg[24][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y31_N3
dffeas \my_reg[20][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][4] .is_wysiwyg = "true";
defparam \my_reg[20][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N2
cycloneive_lcell_comb \Mux27~4 (
// Equation(s):
// \Mux27~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\my_reg[20][4]~q ))) # (!dcifimemload_23 & (\my_reg[16][4]~q ))))

	.dataa(\my_reg[16][4]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[20][4]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~4 .lut_mask = 16'hFC22;
defparam \Mux27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N28
cycloneive_lcell_comb \Mux27~5 (
// Equation(s):
// \Mux27~5_combout  = (dcifimemload_24 & ((\Mux27~4_combout  & (\my_reg[28][4]~q )) # (!\Mux27~4_combout  & ((\my_reg[24][4]~q ))))) # (!dcifimemload_24 & (((\Mux27~4_combout ))))

	.dataa(\my_reg[28][4]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[24][4]~q ),
	.datad(\Mux27~4_combout ),
	.cin(gnd),
	.combout(\Mux27~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~5 .lut_mask = 16'hBBC0;
defparam \Mux27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N0
cycloneive_lcell_comb \my_reg[26][4]~feeder (
// Equation(s):
// \my_reg[26][4]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat29),
	.cin(gnd),
	.combout(\my_reg[26][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[26][4]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[26][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y43_N1
dffeas \my_reg[26][4] (
	.clk(CLK),
	.d(\my_reg[26][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][4] .is_wysiwyg = "true";
defparam \my_reg[26][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N13
dffeas \my_reg[18][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][4] .is_wysiwyg = "true";
defparam \my_reg[18][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N28
cycloneive_lcell_comb \Mux27~2 (
// Equation(s):
// \Mux27~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[22][4]~q )) # (!dcifimemload_23 & ((\my_reg[18][4]~q )))))

	.dataa(\my_reg[22][4]~q ),
	.datab(\my_reg[18][4]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~2 .lut_mask = 16'hFA0C;
defparam \Mux27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N30
cycloneive_lcell_comb \Mux27~3 (
// Equation(s):
// \Mux27~3_combout  = (dcifimemload_24 & ((\Mux27~2_combout  & (\my_reg[30][4]~q )) # (!\Mux27~2_combout  & ((\my_reg[26][4]~q ))))) # (!dcifimemload_24 & (((\Mux27~2_combout ))))

	.dataa(\my_reg[30][4]~q ),
	.datab(\my_reg[26][4]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux27~2_combout ),
	.cin(gnd),
	.combout(\Mux27~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~3 .lut_mask = 16'hAFC0;
defparam \Mux27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N20
cycloneive_lcell_comb \Mux27~6 (
// Equation(s):
// \Mux27~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux27~3_combout ))) # (!dcifimemload_22 & (\Mux27~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux27~5_combout ),
	.datad(\Mux27~3_combout ),
	.cin(gnd),
	.combout(\Mux27~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~6 .lut_mask = 16'hDC98;
defparam \Mux27~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N17
dffeas \my_reg[1][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][4] .is_wysiwyg = "true";
defparam \my_reg[1][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N7
dffeas \my_reg[3][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][4] .is_wysiwyg = "true";
defparam \my_reg[3][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N6
cycloneive_lcell_comb \Mux27~14 (
// Equation(s):
// \Mux27~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][4]~q ))) # (!dcifimemload_22 & (\my_reg[1][4]~q ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[1][4]~q ),
	.datac(\my_reg[3][4]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux27~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~14 .lut_mask = 16'hA088;
defparam \Mux27~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N8
cycloneive_lcell_comb \Mux27~15 (
// Equation(s):
// \Mux27~15_combout  = (\Mux27~14_combout ) # ((\my_reg[2][4]~q  & (dcifimemload_22 & !dcifimemload_21)))

	.dataa(\my_reg[2][4]~q ),
	.datab(\Mux27~14_combout ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux27~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~15 .lut_mask = 16'hCCEC;
defparam \Mux27~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N28
cycloneive_lcell_comb \my_reg[9][4]~feeder (
// Equation(s):
// \my_reg[9][4]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat29),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[9][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[9][4]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[9][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N29
dffeas \my_reg[9][4] (
	.clk(CLK),
	.d(\my_reg[9][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][4] .is_wysiwyg = "true";
defparam \my_reg[9][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N25
dffeas \my_reg[8][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][4] .is_wysiwyg = "true";
defparam \my_reg[8][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N23
dffeas \my_reg[10][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][4] .is_wysiwyg = "true";
defparam \my_reg[10][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N22
cycloneive_lcell_comb \Mux27~12 (
// Equation(s):
// \Mux27~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[10][4]~q ))) # (!dcifimemload_22 & (\my_reg[8][4]~q ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[8][4]~q ),
	.datac(\my_reg[10][4]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux27~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~12 .lut_mask = 16'hFA44;
defparam \Mux27~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N24
cycloneive_lcell_comb \Mux27~13 (
// Equation(s):
// \Mux27~13_combout  = (\Mux27~12_combout  & ((\my_reg[11][4]~q ) # ((!dcifimemload_21)))) # (!\Mux27~12_combout  & (((\my_reg[9][4]~q  & dcifimemload_21))))

	.dataa(\my_reg[11][4]~q ),
	.datab(\my_reg[9][4]~q ),
	.datac(\Mux27~12_combout ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux27~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~13 .lut_mask = 16'hACF0;
defparam \Mux27~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N30
cycloneive_lcell_comb \Mux27~16 (
// Equation(s):
// \Mux27~16_combout  = (dcifimemload_24 & ((dcifimemload_23) # ((\Mux27~13_combout )))) # (!dcifimemload_24 & (!dcifimemload_23 & (\Mux27~15_combout )))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux27~15_combout ),
	.datad(\Mux27~13_combout ),
	.cin(gnd),
	.combout(\Mux27~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~16 .lut_mask = 16'hBA98;
defparam \Mux27~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N19
dffeas \my_reg[15][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][4] .is_wysiwyg = "true";
defparam \my_reg[15][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N8
cycloneive_lcell_comb \my_reg[14][4]~feeder (
// Equation(s):
// \my_reg[14][4]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat29),
	.cin(gnd),
	.combout(\my_reg[14][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[14][4]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[14][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N9
dffeas \my_reg[14][4] (
	.clk(CLK),
	.d(\my_reg[14][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][4] .is_wysiwyg = "true";
defparam \my_reg[14][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N23
dffeas \my_reg[13][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][4] .is_wysiwyg = "true";
defparam \my_reg[13][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N22
cycloneive_lcell_comb \Mux27~17 (
// Equation(s):
// \Mux27~17_combout  = (dcifimemload_21 & (((\my_reg[13][4]~q ) # (dcifimemload_22)))) # (!dcifimemload_21 & (\my_reg[12][4]~q  & ((!dcifimemload_22))))

	.dataa(\my_reg[12][4]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[13][4]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux27~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~17 .lut_mask = 16'hCCE2;
defparam \Mux27~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N30
cycloneive_lcell_comb \Mux27~18 (
// Equation(s):
// \Mux27~18_combout  = (dcifimemload_22 & ((\Mux27~17_combout  & (\my_reg[15][4]~q )) # (!\Mux27~17_combout  & ((\my_reg[14][4]~q ))))) # (!dcifimemload_22 & (((\Mux27~17_combout ))))

	.dataa(\my_reg[15][4]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[14][4]~q ),
	.datad(\Mux27~17_combout ),
	.cin(gnd),
	.combout(\Mux27~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~18 .lut_mask = 16'hBBC0;
defparam \Mux27~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N30
cycloneive_lcell_comb \my_reg[7][4]~feeder (
// Equation(s):
// \my_reg[7][4]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat29),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[7][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[7][4]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[7][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y42_N31
dffeas \my_reg[7][4] (
	.clk(CLK),
	.d(\my_reg[7][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][4] .is_wysiwyg = "true";
defparam \my_reg[7][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N21
dffeas \my_reg[6][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][4] .is_wysiwyg = "true";
defparam \my_reg[6][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N24
cycloneive_lcell_comb \my_reg[4][4]~feeder (
// Equation(s):
// \my_reg[4][4]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat29),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[4][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[4][4]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[4][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y42_N25
dffeas \my_reg[4][4] (
	.clk(CLK),
	.d(\my_reg[4][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][4] .is_wysiwyg = "true";
defparam \my_reg[4][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N3
dffeas \my_reg[5][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][4] .is_wysiwyg = "true";
defparam \my_reg[5][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N2
cycloneive_lcell_comb \Mux27~10 (
// Equation(s):
// \Mux27~10_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\my_reg[5][4]~q ))) # (!dcifimemload_21 & (\my_reg[4][4]~q ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[4][4]~q ),
	.datac(\my_reg[5][4]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux27~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~10 .lut_mask = 16'hFA44;
defparam \Mux27~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N20
cycloneive_lcell_comb \Mux27~11 (
// Equation(s):
// \Mux27~11_combout  = (dcifimemload_22 & ((\Mux27~10_combout  & (\my_reg[7][4]~q )) # (!\Mux27~10_combout  & ((\my_reg[6][4]~q ))))) # (!dcifimemload_22 & (((\Mux27~10_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[7][4]~q ),
	.datac(\my_reg[6][4]~q ),
	.datad(\Mux27~10_combout ),
	.cin(gnd),
	.combout(\Mux27~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~11 .lut_mask = 16'hDDA0;
defparam \Mux27~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N3
dffeas \my_reg[11][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][4] .is_wysiwyg = "true";
defparam \my_reg[11][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N24
cycloneive_lcell_comb \Mux59~0 (
// Equation(s):
// \Mux59~0_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & (\my_reg[10][4]~q )) # (!dcifimemload_17 & ((\my_reg[8][4]~q )))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[10][4]~q ),
	.datac(\my_reg[8][4]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux59~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~0 .lut_mask = 16'hEE50;
defparam \Mux59~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N2
cycloneive_lcell_comb \Mux59~1 (
// Equation(s):
// \Mux59~1_combout  = (dcifimemload_16 & ((\Mux59~0_combout  & ((\my_reg[11][4]~q ))) # (!\Mux59~0_combout  & (\my_reg[9][4]~q )))) # (!dcifimemload_16 & (((\Mux59~0_combout ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[9][4]~q ),
	.datac(\my_reg[11][4]~q ),
	.datad(\Mux59~0_combout ),
	.cin(gnd),
	.combout(\Mux59~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~1 .lut_mask = 16'hF588;
defparam \Mux59~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N25
dffeas \my_reg[12][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][4] .is_wysiwyg = "true";
defparam \my_reg[12][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N24
cycloneive_lcell_comb \Mux59~7 (
// Equation(s):
// \Mux59~7_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\my_reg[13][4]~q )) # (!dcifimemload_16 & ((\my_reg[12][4]~q )))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[13][4]~q ),
	.datac(\my_reg[12][4]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux59~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~7 .lut_mask = 16'hEE50;
defparam \Mux59~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N18
cycloneive_lcell_comb \Mux59~8 (
// Equation(s):
// \Mux59~8_combout  = (dcifimemload_17 & ((\Mux59~7_combout  & ((\my_reg[15][4]~q ))) # (!\Mux59~7_combout  & (\my_reg[14][4]~q )))) # (!dcifimemload_17 & (((\Mux59~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[14][4]~q ),
	.datac(\my_reg[15][4]~q ),
	.datad(\Mux59~7_combout ),
	.cin(gnd),
	.combout(\Mux59~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~8 .lut_mask = 16'hF588;
defparam \Mux59~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N11
dffeas \my_reg[2][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][4] .is_wysiwyg = "true";
defparam \my_reg[2][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N16
cycloneive_lcell_comb \Mux59~4 (
// Equation(s):
// \Mux59~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\my_reg[3][4]~q )) # (!dcifimemload_17 & ((\my_reg[1][4]~q )))))

	.dataa(\my_reg[3][4]~q ),
	.datab(dcifimemload_17),
	.datac(\my_reg[1][4]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux59~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~4 .lut_mask = 16'hB800;
defparam \Mux59~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N10
cycloneive_lcell_comb \Mux59~5 (
// Equation(s):
// \Mux59~5_combout  = (\Mux59~4_combout ) # ((!dcifimemload_16 & (dcifimemload_17 & \my_reg[2][4]~q )))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\my_reg[2][4]~q ),
	.datad(\Mux59~4_combout ),
	.cin(gnd),
	.combout(\Mux59~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~5 .lut_mask = 16'hFF40;
defparam \Mux59~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N20
cycloneive_lcell_comb \Mux59~2 (
// Equation(s):
// \Mux59~2_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\my_reg[5][4]~q )) # (!dcifimemload_16 & ((\my_reg[4][4]~q )))))

	.dataa(\my_reg[5][4]~q ),
	.datab(\my_reg[4][4]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux59~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~2 .lut_mask = 16'hFA0C;
defparam \Mux59~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N22
cycloneive_lcell_comb \Mux59~3 (
// Equation(s):
// \Mux59~3_combout  = (dcifimemload_17 & ((\Mux59~2_combout  & (\my_reg[7][4]~q )) # (!\Mux59~2_combout  & ((\my_reg[6][4]~q ))))) # (!dcifimemload_17 & (((\Mux59~2_combout ))))

	.dataa(\my_reg[7][4]~q ),
	.datab(\my_reg[6][4]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux59~2_combout ),
	.cin(gnd),
	.combout(\Mux59~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~3 .lut_mask = 16'hAFC0;
defparam \Mux59~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N0
cycloneive_lcell_comb \Mux59~6 (
// Equation(s):
// \Mux59~6_combout  = (dcifimemload_18 & ((dcifimemload_19) # ((\Mux59~3_combout )))) # (!dcifimemload_18 & (!dcifimemload_19 & (\Mux59~5_combout )))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux59~5_combout ),
	.datad(\Mux59~3_combout ),
	.cin(gnd),
	.combout(\Mux59~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~6 .lut_mask = 16'hBA98;
defparam \Mux59~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N2
cycloneive_lcell_comb \Mux59~17 (
// Equation(s):
// \Mux59~17_combout  = (dcifimemload_18 & (((\my_reg[23][4]~q ) # (dcifimemload_19)))) # (!dcifimemload_18 & (\my_reg[19][4]~q  & ((!dcifimemload_19))))

	.dataa(\my_reg[19][4]~q ),
	.datab(\my_reg[23][4]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux59~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~17 .lut_mask = 16'hF0CA;
defparam \Mux59~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N4
cycloneive_lcell_comb \Mux59~18 (
// Equation(s):
// \Mux59~18_combout  = (dcifimemload_19 & ((\Mux59~17_combout  & (\my_reg[31][4]~q )) # (!\Mux59~17_combout  & ((\my_reg[27][4]~q ))))) # (!dcifimemload_19 & (((\Mux59~17_combout ))))

	.dataa(\my_reg[31][4]~q ),
	.datab(\my_reg[27][4]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux59~17_combout ),
	.cin(gnd),
	.combout(\Mux59~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~18 .lut_mask = 16'hAFC0;
defparam \Mux59~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N23
dffeas \my_reg[28][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][4] .is_wysiwyg = "true";
defparam \my_reg[28][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N17
dffeas \my_reg[16][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][4] .is_wysiwyg = "true";
defparam \my_reg[16][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N16
cycloneive_lcell_comb \Mux59~14 (
// Equation(s):
// \Mux59~14_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\my_reg[24][4]~q )) # (!dcifimemload_19 & ((\my_reg[16][4]~q )))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[24][4]~q ),
	.datac(\my_reg[16][4]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux59~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~14 .lut_mask = 16'hEE50;
defparam \Mux59~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N22
cycloneive_lcell_comb \Mux59~15 (
// Equation(s):
// \Mux59~15_combout  = (dcifimemload_18 & ((\Mux59~14_combout  & ((\my_reg[28][4]~q ))) # (!\Mux59~14_combout  & (\my_reg[20][4]~q )))) # (!dcifimemload_18 & (((\Mux59~14_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[20][4]~q ),
	.datac(\my_reg[28][4]~q ),
	.datad(\Mux59~14_combout ),
	.cin(gnd),
	.combout(\Mux59~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~15 .lut_mask = 16'hF588;
defparam \Mux59~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N6
cycloneive_lcell_comb \my_reg[22][4]~feeder (
// Equation(s):
// \my_reg[22][4]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat29),
	.cin(gnd),
	.combout(\my_reg[22][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[22][4]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[22][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y43_N7
dffeas \my_reg[22][4] (
	.clk(CLK),
	.d(\my_reg[22][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][4] .is_wysiwyg = "true";
defparam \my_reg[22][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N31
dffeas \my_reg[30][4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][4] .is_wysiwyg = "true";
defparam \my_reg[30][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N12
cycloneive_lcell_comb \Mux59~12 (
// Equation(s):
// \Mux59~12_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\my_reg[26][4]~q )) # (!dcifimemload_19 & ((\my_reg[18][4]~q )))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[26][4]~q ),
	.datac(\my_reg[18][4]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux59~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~12 .lut_mask = 16'hEE50;
defparam \Mux59~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N30
cycloneive_lcell_comb \Mux59~13 (
// Equation(s):
// \Mux59~13_combout  = (dcifimemload_18 & ((\Mux59~12_combout  & ((\my_reg[30][4]~q ))) # (!\Mux59~12_combout  & (\my_reg[22][4]~q )))) # (!dcifimemload_18 & (((\Mux59~12_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[22][4]~q ),
	.datac(\my_reg[30][4]~q ),
	.datad(\Mux59~12_combout ),
	.cin(gnd),
	.combout(\Mux59~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~13 .lut_mask = 16'hF588;
defparam \Mux59~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N26
cycloneive_lcell_comb \Mux59~16 (
// Equation(s):
// \Mux59~16_combout  = (dcifimemload_16 & (((dcifimemload_17)))) # (!dcifimemload_16 & ((dcifimemload_17 & ((\Mux59~13_combout ))) # (!dcifimemload_17 & (\Mux59~15_combout ))))

	.dataa(\Mux59~15_combout ),
	.datab(dcifimemload_16),
	.datac(\Mux59~13_combout ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux59~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~16 .lut_mask = 16'hFC22;
defparam \Mux59~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N28
cycloneive_lcell_comb \my_reg[17][4]~feeder (
// Equation(s):
// \my_reg[17][4]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat29),
	.cin(gnd),
	.combout(\my_reg[17][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[17][4]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[17][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y40_N29
dffeas \my_reg[17][4] (
	.clk(CLK),
	.d(\my_reg[17][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][4] .is_wysiwyg = "true";
defparam \my_reg[17][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N30
cycloneive_lcell_comb \Mux59~10 (
// Equation(s):
// \Mux59~10_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\my_reg[21][4]~q )) # (!dcifimemload_18 & ((\my_reg[17][4]~q )))))

	.dataa(\my_reg[21][4]~q ),
	.datab(\my_reg[17][4]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux59~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~10 .lut_mask = 16'hFA0C;
defparam \Mux59~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N24
cycloneive_lcell_comb \Mux59~11 (
// Equation(s):
// \Mux59~11_combout  = (dcifimemload_19 & ((\Mux59~10_combout  & ((\my_reg[29][4]~q ))) # (!\Mux59~10_combout  & (\my_reg[25][4]~q )))) # (!dcifimemload_19 & (((\Mux59~10_combout ))))

	.dataa(\my_reg[25][4]~q ),
	.datab(\my_reg[29][4]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux59~10_combout ),
	.cin(gnd),
	.combout(\Mux59~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~11 .lut_mask = 16'hCFA0;
defparam \Mux59~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N22
cycloneive_lcell_comb \my_reg[14][3]~feeder (
// Equation(s):
// \my_reg[14][3]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat30),
	.cin(gnd),
	.combout(\my_reg[14][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[14][3]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[14][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N23
dffeas \my_reg[14][3] (
	.clk(CLK),
	.d(\my_reg[14][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][3] .is_wysiwyg = "true";
defparam \my_reg[14][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N12
cycloneive_lcell_comb \my_reg[12][3]~feeder (
// Equation(s):
// \my_reg[12][3]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat30),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[12][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[12][3]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[12][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N13
dffeas \my_reg[12][3] (
	.clk(CLK),
	.d(\my_reg[12][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][3] .is_wysiwyg = "true";
defparam \my_reg[12][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N13
dffeas \my_reg[13][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][3] .is_wysiwyg = "true";
defparam \my_reg[13][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N12
cycloneive_lcell_comb \Mux28~17 (
// Equation(s):
// \Mux28~17_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\my_reg[13][3]~q ))) # (!dcifimemload_21 & (\my_reg[12][3]~q ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[12][3]~q ),
	.datac(\my_reg[13][3]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux28~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~17 .lut_mask = 16'hFA44;
defparam \Mux28~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N27
dffeas \my_reg[15][3] (
	.clk(CLK),
	.d(wdat30),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][3] .is_wysiwyg = "true";
defparam \my_reg[15][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N8
cycloneive_lcell_comb \Mux28~18 (
// Equation(s):
// \Mux28~18_combout  = (dcifimemload_22 & ((\Mux28~17_combout  & ((\my_reg[15][3]~q ))) # (!\Mux28~17_combout  & (\my_reg[14][3]~q )))) # (!dcifimemload_22 & (((\Mux28~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[14][3]~q ),
	.datac(\Mux28~17_combout ),
	.datad(\my_reg[15][3]~q ),
	.cin(gnd),
	.combout(\Mux28~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~18 .lut_mask = 16'hF858;
defparam \Mux28~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N31
dffeas \my_reg[7][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][3] .is_wysiwyg = "true";
defparam \my_reg[7][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N17
dffeas \my_reg[4][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][3] .is_wysiwyg = "true";
defparam \my_reg[4][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N16
cycloneive_lcell_comb \Mux28~12 (
// Equation(s):
// \Mux28~12_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & (\my_reg[5][3]~q )) # (!dcifimemload_21 & ((\my_reg[4][3]~q )))))

	.dataa(\my_reg[5][3]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[4][3]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux28~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~12 .lut_mask = 16'hEE30;
defparam \Mux28~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N30
cycloneive_lcell_comb \Mux28~13 (
// Equation(s):
// \Mux28~13_combout  = (dcifimemload_22 & ((\Mux28~12_combout  & ((\my_reg[7][3]~q ))) # (!\Mux28~12_combout  & (\my_reg[6][3]~q )))) # (!dcifimemload_22 & (((\Mux28~12_combout ))))

	.dataa(\my_reg[6][3]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[7][3]~q ),
	.datad(\Mux28~12_combout ),
	.cin(gnd),
	.combout(\Mux28~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~13 .lut_mask = 16'hF388;
defparam \Mux28~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N15
dffeas \my_reg[2][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][3] .is_wysiwyg = "true";
defparam \my_reg[2][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N28
cycloneive_lcell_comb \my_reg[3][3]~feeder (
// Equation(s):
// \my_reg[3][3]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat30),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[3][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[3][3]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[3][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y37_N29
dffeas \my_reg[3][3] (
	.clk(CLK),
	.d(\my_reg[3][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][3] .is_wysiwyg = "true";
defparam \my_reg[3][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N10
cycloneive_lcell_comb \Mux28~14 (
// Equation(s):
// \Mux28~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][3]~q ))) # (!dcifimemload_22 & (\my_reg[1][3]~q ))))

	.dataa(\my_reg[1][3]~q ),
	.datab(\my_reg[3][3]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux28~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~14 .lut_mask = 16'hCA00;
defparam \Mux28~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N12
cycloneive_lcell_comb \Mux28~15 (
// Equation(s):
// \Mux28~15_combout  = (\Mux28~14_combout ) # ((dcifimemload_22 & (\my_reg[2][3]~q  & !dcifimemload_21)))

	.dataa(dcifimemload_22),
	.datab(\my_reg[2][3]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux28~14_combout ),
	.cin(gnd),
	.combout(\Mux28~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~15 .lut_mask = 16'hFF08;
defparam \Mux28~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N30
cycloneive_lcell_comb \Mux28~16 (
// Equation(s):
// \Mux28~16_combout  = (dcifimemload_24 & (dcifimemload_23)) # (!dcifimemload_24 & ((dcifimemload_23 & (\Mux28~13_combout )) # (!dcifimemload_23 & ((\Mux28~15_combout )))))

	.dataa(dcifimemload_24),
	.datab(dcifimemload_23),
	.datac(\Mux28~13_combout ),
	.datad(\Mux28~15_combout ),
	.cin(gnd),
	.combout(\Mux28~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~16 .lut_mask = 16'hD9C8;
defparam \Mux28~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N19
dffeas \my_reg[11][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][3] .is_wysiwyg = "true";
defparam \my_reg[11][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N29
dffeas \my_reg[9][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][3] .is_wysiwyg = "true";
defparam \my_reg[9][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N29
dffeas \my_reg[8][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][3] .is_wysiwyg = "true";
defparam \my_reg[8][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N11
dffeas \my_reg[10][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[10][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[10][3] .is_wysiwyg = "true";
defparam \my_reg[10][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N10
cycloneive_lcell_comb \Mux28~10 (
// Equation(s):
// \Mux28~10_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[10][3]~q ))) # (!dcifimemload_22 & (\my_reg[8][3]~q ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[8][3]~q ),
	.datac(\my_reg[10][3]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux28~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~10 .lut_mask = 16'hFA44;
defparam \Mux28~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N28
cycloneive_lcell_comb \Mux28~11 (
// Equation(s):
// \Mux28~11_combout  = (dcifimemload_21 & ((\Mux28~10_combout  & (\my_reg[11][3]~q )) # (!\Mux28~10_combout  & ((\my_reg[9][3]~q ))))) # (!dcifimemload_21 & (((\Mux28~10_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[11][3]~q ),
	.datac(\my_reg[9][3]~q ),
	.datad(\Mux28~10_combout ),
	.cin(gnd),
	.combout(\Mux28~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~11 .lut_mask = 16'hDDA0;
defparam \Mux28~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N26
cycloneive_lcell_comb \Mux28~19 (
// Equation(s):
// \Mux28~19_combout  = (dcifimemload_24 & ((\Mux28~16_combout  & (\Mux28~18_combout )) # (!\Mux28~16_combout  & ((\Mux28~11_combout ))))) # (!dcifimemload_24 & (((\Mux28~16_combout ))))

	.dataa(dcifimemload_24),
	.datab(\Mux28~18_combout ),
	.datac(\Mux28~16_combout ),
	.datad(\Mux28~11_combout ),
	.cin(gnd),
	.combout(\Mux28~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~19 .lut_mask = 16'hDAD0;
defparam \Mux28~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N15
dffeas \my_reg[29][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][3] .is_wysiwyg = "true";
defparam \my_reg[29][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N13
dffeas \my_reg[17][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][3] .is_wysiwyg = "true";
defparam \my_reg[17][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N12
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[21][3]~q )) # (!dcifimemload_23 & ((\my_reg[17][3]~q )))))

	.dataa(\my_reg[21][3]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[17][3]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'hEE30;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N14
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (dcifimemload_24 & ((\Mux28~0_combout  & ((\my_reg[29][3]~q ))) # (!\Mux28~0_combout  & (\my_reg[25][3]~q )))) # (!dcifimemload_24 & (((\Mux28~0_combout ))))

	.dataa(\my_reg[25][3]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[29][3]~q ),
	.datad(\Mux28~0_combout ),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hF388;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N14
cycloneive_lcell_comb \my_reg[31][3]~feeder (
// Equation(s):
// \my_reg[31][3]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat30),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[31][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[31][3]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[31][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N15
dffeas \my_reg[31][3] (
	.clk(CLK),
	.d(\my_reg[31][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][3] .is_wysiwyg = "true";
defparam \my_reg[31][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y35_N7
dffeas \my_reg[27][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][3] .is_wysiwyg = "true";
defparam \my_reg[27][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N23
dffeas \my_reg[23][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][3] .is_wysiwyg = "true";
defparam \my_reg[23][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N22
cycloneive_lcell_comb \Mux28~7 (
// Equation(s):
// \Mux28~7_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & ((\my_reg[23][3]~q ))) # (!dcifimemload_23 & (\my_reg[19][3]~q ))))

	.dataa(\my_reg[19][3]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[23][3]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux28~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~7 .lut_mask = 16'hFC22;
defparam \Mux28~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N6
cycloneive_lcell_comb \Mux28~8 (
// Equation(s):
// \Mux28~8_combout  = (dcifimemload_24 & ((\Mux28~7_combout  & (\my_reg[31][3]~q )) # (!\Mux28~7_combout  & ((\my_reg[27][3]~q ))))) # (!dcifimemload_24 & (((\Mux28~7_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[31][3]~q ),
	.datac(\my_reg[27][3]~q ),
	.datad(\Mux28~7_combout ),
	.cin(gnd),
	.combout(\Mux28~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~8 .lut_mask = 16'hDDA0;
defparam \Mux28~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N1
dffeas \my_reg[30][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][3] .is_wysiwyg = "true";
defparam \my_reg[30][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N14
cycloneive_lcell_comb \my_reg[18][3]~feeder (
// Equation(s):
// \my_reg[18][3]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat30),
	.cin(gnd),
	.combout(\my_reg[18][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[18][3]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[18][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y30_N15
dffeas \my_reg[18][3] (
	.clk(CLK),
	.d(\my_reg[18][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][3] .is_wysiwyg = "true";
defparam \my_reg[18][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N8
cycloneive_lcell_comb \Mux28~2 (
// Equation(s):
// \Mux28~2_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[26][3]~q )) # (!dcifimemload_24 & ((\my_reg[18][3]~q )))))

	.dataa(\my_reg[26][3]~q ),
	.datab(\my_reg[18][3]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~2 .lut_mask = 16'hFA0C;
defparam \Mux28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N0
cycloneive_lcell_comb \Mux28~3 (
// Equation(s):
// \Mux28~3_combout  = (dcifimemload_23 & ((\Mux28~2_combout  & ((\my_reg[30][3]~q ))) # (!\Mux28~2_combout  & (\my_reg[22][3]~q )))) # (!dcifimemload_23 & (((\Mux28~2_combout ))))

	.dataa(\my_reg[22][3]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[30][3]~q ),
	.datad(\Mux28~2_combout ),
	.cin(gnd),
	.combout(\Mux28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~3 .lut_mask = 16'hF388;
defparam \Mux28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N28
cycloneive_lcell_comb \Mux28~6 (
// Equation(s):
// \Mux28~6_combout  = (dcifimemload_22 & (((dcifimemload_21) # (\Mux28~3_combout )))) # (!dcifimemload_22 & (\Mux28~5_combout  & (!dcifimemload_21)))

	.dataa(\Mux28~5_combout ),
	.datab(dcifimemload_22),
	.datac(dcifimemload_21),
	.datad(\Mux28~3_combout ),
	.cin(gnd),
	.combout(\Mux28~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~6 .lut_mask = 16'hCEC2;
defparam \Mux28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N2
cycloneive_lcell_comb \Mux28~9 (
// Equation(s):
// \Mux28~9_combout  = (dcifimemload_21 & ((\Mux28~6_combout  & ((\Mux28~8_combout ))) # (!\Mux28~6_combout  & (\Mux28~1_combout )))) # (!dcifimemload_21 & (((\Mux28~6_combout ))))

	.dataa(dcifimemload_21),
	.datab(\Mux28~1_combout ),
	.datac(\Mux28~8_combout ),
	.datad(\Mux28~6_combout ),
	.cin(gnd),
	.combout(\Mux28~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~9 .lut_mask = 16'hF588;
defparam \Mux28~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N12
cycloneive_lcell_comb \my_reg[19][3]~feeder (
// Equation(s):
// \my_reg[19][3]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat30),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[19][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[19][3]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[19][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y34_N13
dffeas \my_reg[19][3] (
	.clk(CLK),
	.d(\my_reg[19][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][3] .is_wysiwyg = "true";
defparam \my_reg[19][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N16
cycloneive_lcell_comb \Mux60~7 (
// Equation(s):
// \Mux60~7_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\my_reg[27][3]~q )) # (!dcifimemload_19 & ((\my_reg[19][3]~q )))))

	.dataa(\my_reg[27][3]~q ),
	.datab(\my_reg[19][3]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux60~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~7 .lut_mask = 16'hFA0C;
defparam \Mux60~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N18
cycloneive_lcell_comb \Mux60~8 (
// Equation(s):
// \Mux60~8_combout  = (dcifimemload_18 & ((\Mux60~7_combout  & (\my_reg[31][3]~q )) # (!\Mux60~7_combout  & ((\my_reg[23][3]~q ))))) # (!dcifimemload_18 & (((\Mux60~7_combout ))))

	.dataa(\my_reg[31][3]~q ),
	.datab(\my_reg[23][3]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux60~7_combout ),
	.cin(gnd),
	.combout(\Mux60~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~8 .lut_mask = 16'hAFC0;
defparam \Mux60~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N14
cycloneive_lcell_comb \my_reg[21][3]~feeder (
// Equation(s):
// \my_reg[21][3]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat30),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[21][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[21][3]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[21][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y35_N15
dffeas \my_reg[21][3] (
	.clk(CLK),
	.d(\my_reg[21][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][3] .is_wysiwyg = "true";
defparam \my_reg[21][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N12
cycloneive_lcell_comb \my_reg[25][3]~feeder (
// Equation(s):
// \my_reg[25][3]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat30),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[25][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[25][3]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[25][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y35_N13
dffeas \my_reg[25][3] (
	.clk(CLK),
	.d(\my_reg[25][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][3] .is_wysiwyg = "true";
defparam \my_reg[25][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N0
cycloneive_lcell_comb \Mux60~0 (
// Equation(s):
// \Mux60~0_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & ((\my_reg[25][3]~q ))) # (!dcifimemload_19 & (\my_reg[17][3]~q ))))

	.dataa(\my_reg[17][3]~q ),
	.datab(\my_reg[25][3]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux60~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~0 .lut_mask = 16'hFC0A;
defparam \Mux60~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N6
cycloneive_lcell_comb \Mux60~1 (
// Equation(s):
// \Mux60~1_combout  = (dcifimemload_18 & ((\Mux60~0_combout  & (\my_reg[29][3]~q )) # (!\Mux60~0_combout  & ((\my_reg[21][3]~q ))))) # (!dcifimemload_18 & (((\Mux60~0_combout ))))

	.dataa(\my_reg[29][3]~q ),
	.datab(\my_reg[21][3]~q ),
	.datac(dcifimemload_18),
	.datad(\Mux60~0_combout ),
	.cin(gnd),
	.combout(\Mux60~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~1 .lut_mask = 16'hAFC0;
defparam \Mux60~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N20
cycloneive_lcell_comb \my_reg[26][3]~feeder (
// Equation(s):
// \my_reg[26][3]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat30),
	.cin(gnd),
	.combout(\my_reg[26][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[26][3]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[26][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y30_N21
dffeas \my_reg[26][3] (
	.clk(CLK),
	.d(\my_reg[26][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][3] .is_wysiwyg = "true";
defparam \my_reg[26][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N19
dffeas \my_reg[22][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][3] .is_wysiwyg = "true";
defparam \my_reg[22][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N18
cycloneive_lcell_comb \Mux60~2 (
// Equation(s):
// \Mux60~2_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[22][3]~q ))) # (!dcifimemload_18 & (\my_reg[18][3]~q ))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[18][3]~q ),
	.datac(\my_reg[22][3]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux60~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~2 .lut_mask = 16'hFA44;
defparam \Mux60~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y30_N10
cycloneive_lcell_comb \Mux60~3 (
// Equation(s):
// \Mux60~3_combout  = (\Mux60~2_combout  & ((\my_reg[30][3]~q ) # ((!dcifimemload_19)))) # (!\Mux60~2_combout  & (((\my_reg[26][3]~q  & dcifimemload_19))))

	.dataa(\my_reg[30][3]~q ),
	.datab(\my_reg[26][3]~q ),
	.datac(\Mux60~2_combout ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux60~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~3 .lut_mask = 16'hACF0;
defparam \Mux60~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N24
cycloneive_lcell_comb \my_reg[28][3]~feeder (
// Equation(s):
// \my_reg[28][3]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat30),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[28][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[28][3]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[28][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N25
dffeas \my_reg[28][3] (
	.clk(CLK),
	.d(\my_reg[28][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][3] .is_wysiwyg = "true";
defparam \my_reg[28][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N28
cycloneive_lcell_comb \my_reg[20][3]~feeder (
// Equation(s):
// \my_reg[20][3]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat30),
	.cin(gnd),
	.combout(\my_reg[20][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[20][3]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[20][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y29_N29
dffeas \my_reg[20][3] (
	.clk(CLK),
	.d(\my_reg[20][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[20][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[20][3] .is_wysiwyg = "true";
defparam \my_reg[20][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N20
cycloneive_lcell_comb \Mux60~4 (
// Equation(s):
// \Mux60~4_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[20][3]~q ))) # (!dcifimemload_18 & (\my_reg[16][3]~q ))))

	.dataa(\my_reg[16][3]~q ),
	.datab(\my_reg[20][3]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux60~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~4 .lut_mask = 16'hFC0A;
defparam \Mux60~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N30
cycloneive_lcell_comb \Mux60~5 (
// Equation(s):
// \Mux60~5_combout  = (dcifimemload_19 & ((\Mux60~4_combout  & ((\my_reg[28][3]~q ))) # (!\Mux60~4_combout  & (\my_reg[24][3]~q )))) # (!dcifimemload_19 & (((\Mux60~4_combout ))))

	.dataa(\my_reg[24][3]~q ),
	.datab(\my_reg[28][3]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux60~4_combout ),
	.cin(gnd),
	.combout(\Mux60~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~5 .lut_mask = 16'hCFA0;
defparam \Mux60~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N20
cycloneive_lcell_comb \Mux60~6 (
// Equation(s):
// \Mux60~6_combout  = (dcifimemload_16 & (dcifimemload_17)) # (!dcifimemload_16 & ((dcifimemload_17 & (\Mux60~3_combout )) # (!dcifimemload_17 & ((\Mux60~5_combout )))))

	.dataa(dcifimemload_16),
	.datab(dcifimemload_17),
	.datac(\Mux60~3_combout ),
	.datad(\Mux60~5_combout ),
	.cin(gnd),
	.combout(\Mux60~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~6 .lut_mask = 16'hD9C8;
defparam \Mux60~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y32_N13
dffeas \my_reg[6][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][3] .is_wysiwyg = "true";
defparam \my_reg[6][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y32_N7
dffeas \my_reg[5][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][3] .is_wysiwyg = "true";
defparam \my_reg[5][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N6
cycloneive_lcell_comb \Mux60~10 (
// Equation(s):
// \Mux60~10_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][3]~q ))) # (!dcifimemload_16 & (\my_reg[4][3]~q ))))

	.dataa(\my_reg[4][3]~q ),
	.datab(dcifimemload_17),
	.datac(\my_reg[5][3]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux60~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~10 .lut_mask = 16'hFC22;
defparam \Mux60~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N12
cycloneive_lcell_comb \Mux60~11 (
// Equation(s):
// \Mux60~11_combout  = (dcifimemload_17 & ((\Mux60~10_combout  & (\my_reg[7][3]~q )) # (!\Mux60~10_combout  & ((\my_reg[6][3]~q ))))) # (!dcifimemload_17 & (((\Mux60~10_combout ))))

	.dataa(\my_reg[7][3]~q ),
	.datab(dcifimemload_17),
	.datac(\my_reg[6][3]~q ),
	.datad(\Mux60~10_combout ),
	.cin(gnd),
	.combout(\Mux60~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~11 .lut_mask = 16'hBBC0;
defparam \Mux60~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N16
cycloneive_lcell_comb \Mux60~17 (
// Equation(s):
// \Mux60~17_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & (\my_reg[13][3]~q )) # (!dcifimemload_16 & ((\my_reg[12][3]~q )))))

	.dataa(\my_reg[13][3]~q ),
	.datab(\my_reg[12][3]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux60~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~17 .lut_mask = 16'hFA0C;
defparam \Mux60~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N2
cycloneive_lcell_comb \Mux60~18 (
// Equation(s):
// \Mux60~18_combout  = (dcifimemload_17 & ((\Mux60~17_combout  & ((\my_reg[15][3]~q ))) # (!\Mux60~17_combout  & (\my_reg[14][3]~q )))) # (!dcifimemload_17 & (((\Mux60~17_combout ))))

	.dataa(\my_reg[14][3]~q ),
	.datab(\my_reg[15][3]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux60~17_combout ),
	.cin(gnd),
	.combout(\Mux60~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~18 .lut_mask = 16'hCFA0;
defparam \Mux60~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N21
dffeas \my_reg[1][3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][3] .is_wysiwyg = "true";
defparam \my_reg[1][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N20
cycloneive_lcell_comb \Mux60~14 (
// Equation(s):
// \Mux60~14_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\my_reg[3][3]~q )) # (!dcifimemload_17 & ((\my_reg[1][3]~q )))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[3][3]~q ),
	.datac(\my_reg[1][3]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux60~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~14 .lut_mask = 16'hD800;
defparam \Mux60~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N14
cycloneive_lcell_comb \Mux60~15 (
// Equation(s):
// \Mux60~15_combout  = (\Mux60~14_combout ) # ((dcifimemload_17 & (\my_reg[2][3]~q  & !dcifimemload_16)))

	.dataa(dcifimemload_17),
	.datab(\Mux60~14_combout ),
	.datac(\my_reg[2][3]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux60~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~15 .lut_mask = 16'hCCEC;
defparam \Mux60~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N28
cycloneive_lcell_comb \Mux60~12 (
// Equation(s):
// \Mux60~12_combout  = (dcifimemload_17 & ((\my_reg[10][3]~q ) # ((dcifimemload_16)))) # (!dcifimemload_17 & (((\my_reg[8][3]~q  & !dcifimemload_16))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[10][3]~q ),
	.datac(\my_reg[8][3]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux60~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~12 .lut_mask = 16'hAAD8;
defparam \Mux60~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N18
cycloneive_lcell_comb \Mux60~13 (
// Equation(s):
// \Mux60~13_combout  = (dcifimemload_16 & ((\Mux60~12_combout  & ((\my_reg[11][3]~q ))) # (!\Mux60~12_combout  & (\my_reg[9][3]~q )))) # (!dcifimemload_16 & (((\Mux60~12_combout ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[9][3]~q ),
	.datac(\my_reg[11][3]~q ),
	.datad(\Mux60~12_combout ),
	.cin(gnd),
	.combout(\Mux60~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~13 .lut_mask = 16'hF588;
defparam \Mux60~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N12
cycloneive_lcell_comb \Mux60~16 (
// Equation(s):
// \Mux60~16_combout  = (dcifimemload_18 & (dcifimemload_19)) # (!dcifimemload_18 & ((dcifimemload_19 & ((\Mux60~13_combout ))) # (!dcifimemload_19 & (\Mux60~15_combout ))))

	.dataa(dcifimemload_18),
	.datab(dcifimemload_19),
	.datac(\Mux60~15_combout ),
	.datad(\Mux60~13_combout ),
	.cin(gnd),
	.combout(\Mux60~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~16 .lut_mask = 16'hDC98;
defparam \Mux60~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N10
cycloneive_lcell_comb \my_reg[31][2]~feeder (
// Equation(s):
// \my_reg[31][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat31),
	.cin(gnd),
	.combout(\my_reg[31][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[31][2]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[31][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N11
dffeas \my_reg[31][2] (
	.clk(CLK),
	.d(\my_reg[31][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[31][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[31][2] .is_wysiwyg = "true";
defparam \my_reg[31][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N24
cycloneive_lcell_comb \my_reg[23][2]~feeder (
// Equation(s):
// \my_reg[23][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat31),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[23][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[23][2]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[23][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N25
dffeas \my_reg[23][2] (
	.clk(CLK),
	.d(\my_reg[23][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[23][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[23][2] .is_wysiwyg = "true";
defparam \my_reg[23][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N24
cycloneive_lcell_comb \my_reg[19][2]~feeder (
// Equation(s):
// \my_reg[19][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat31),
	.cin(gnd),
	.combout(\my_reg[19][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[19][2]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[19][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N25
dffeas \my_reg[19][2] (
	.clk(CLK),
	.d(\my_reg[19][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][2] .is_wysiwyg = "true";
defparam \my_reg[19][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N0
cycloneive_lcell_comb \Mux29~7 (
// Equation(s):
// \Mux29~7_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[27][2]~q )) # (!dcifimemload_24 & ((\my_reg[19][2]~q )))))

	.dataa(\my_reg[27][2]~q ),
	.datab(\my_reg[19][2]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux29~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~7 .lut_mask = 16'hFA0C;
defparam \Mux29~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N18
cycloneive_lcell_comb \Mux29~8 (
// Equation(s):
// \Mux29~8_combout  = (dcifimemload_23 & ((\Mux29~7_combout  & (\my_reg[31][2]~q )) # (!\Mux29~7_combout  & ((\my_reg[23][2]~q ))))) # (!dcifimemload_23 & (((\Mux29~7_combout ))))

	.dataa(\my_reg[31][2]~q ),
	.datab(\my_reg[23][2]~q ),
	.datac(dcifimemload_23),
	.datad(\Mux29~7_combout ),
	.cin(gnd),
	.combout(\Mux29~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~8 .lut_mask = 16'hAFC0;
defparam \Mux29~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y31_N5
dffeas \my_reg[21][2] (
	.clk(CLK),
	.d(wdat31),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[21][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[21][2] .is_wysiwyg = "true";
defparam \my_reg[21][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N15
dffeas \my_reg[25][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[25][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[25][2] .is_wysiwyg = "true";
defparam \my_reg[25][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N14
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (dcifimemload_24 & (((\my_reg[25][2]~q ) # (dcifimemload_23)))) # (!dcifimemload_24 & (\my_reg[17][2]~q  & ((!dcifimemload_23))))

	.dataa(\my_reg[17][2]~q ),
	.datab(dcifimemload_24),
	.datac(\my_reg[25][2]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hCCE2;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N0
cycloneive_lcell_comb \my_reg[29][2]~feeder (
// Equation(s):
// \my_reg[29][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat31),
	.cin(gnd),
	.combout(\my_reg[29][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[29][2]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[29][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N1
dffeas \my_reg[29][2] (
	.clk(CLK),
	.d(\my_reg[29][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[29][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[29][2] .is_wysiwyg = "true";
defparam \my_reg[29][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N22
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// \Mux29~1_combout  = (\Mux29~0_combout  & (((\my_reg[29][2]~q ) # (!dcifimemload_23)))) # (!\Mux29~0_combout  & (\my_reg[21][2]~q  & ((dcifimemload_23))))

	.dataa(\my_reg[21][2]~q ),
	.datab(\Mux29~0_combout ),
	.datac(\my_reg[29][2]~q ),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hE2CC;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N8
cycloneive_lcell_comb \my_reg[24][2]~feeder (
// Equation(s):
// \my_reg[24][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat31),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[24][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[24][2]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[24][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y31_N9
dffeas \my_reg[24][2] (
	.clk(CLK),
	.d(\my_reg[24][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[24][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[24][2] .is_wysiwyg = "true";
defparam \my_reg[24][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N21
dffeas \my_reg[16][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[16][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[16][2] .is_wysiwyg = "true";
defparam \my_reg[16][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N20
cycloneive_lcell_comb \Mux29~4 (
// Equation(s):
// \Mux29~4_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[20][2]~q )) # (!dcifimemload_23 & ((\my_reg[16][2]~q )))))

	.dataa(\my_reg[20][2]~q ),
	.datab(\my_reg[16][2]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~4 .lut_mask = 16'hFA0C;
defparam \Mux29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N22
cycloneive_lcell_comb \Mux29~5 (
// Equation(s):
// \Mux29~5_combout  = (dcifimemload_24 & ((\Mux29~4_combout  & (\my_reg[28][2]~q )) # (!\Mux29~4_combout  & ((\my_reg[24][2]~q ))))) # (!dcifimemload_24 & (((\Mux29~4_combout ))))

	.dataa(\my_reg[28][2]~q ),
	.datab(\my_reg[24][2]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux29~4_combout ),
	.cin(gnd),
	.combout(\Mux29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~5 .lut_mask = 16'hAFC0;
defparam \Mux29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N27
dffeas \my_reg[30][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[30][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[30][2] .is_wysiwyg = "true";
defparam \my_reg[30][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N17
dffeas \my_reg[18][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[18][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[18][2] .is_wysiwyg = "true";
defparam \my_reg[18][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N12
cycloneive_lcell_comb \Mux29~2 (
// Equation(s):
// \Mux29~2_combout  = (dcifimemload_24 & (((dcifimemload_23)))) # (!dcifimemload_24 & ((dcifimemload_23 & (\my_reg[22][2]~q )) # (!dcifimemload_23 & ((\my_reg[18][2]~q )))))

	.dataa(\my_reg[22][2]~q ),
	.datab(\my_reg[18][2]~q ),
	.datac(dcifimemload_24),
	.datad(dcifimemload_23),
	.cin(gnd),
	.combout(\Mux29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~2 .lut_mask = 16'hFA0C;
defparam \Mux29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N2
cycloneive_lcell_comb \Mux29~3 (
// Equation(s):
// \Mux29~3_combout  = (dcifimemload_24 & ((\Mux29~2_combout  & ((\my_reg[30][2]~q ))) # (!\Mux29~2_combout  & (\my_reg[26][2]~q )))) # (!dcifimemload_24 & (((\Mux29~2_combout ))))

	.dataa(\my_reg[26][2]~q ),
	.datab(\my_reg[30][2]~q ),
	.datac(dcifimemload_24),
	.datad(\Mux29~2_combout ),
	.cin(gnd),
	.combout(\Mux29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~3 .lut_mask = 16'hCFA0;
defparam \Mux29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N24
cycloneive_lcell_comb \Mux29~6 (
// Equation(s):
// \Mux29~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & ((\Mux29~3_combout ))) # (!dcifimemload_22 & (\Mux29~5_combout ))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux29~5_combout ),
	.datad(\Mux29~3_combout ),
	.cin(gnd),
	.combout(\Mux29~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~6 .lut_mask = 16'hDC98;
defparam \Mux29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N24
cycloneive_lcell_comb \my_reg[14][2]~feeder (
// Equation(s):
// \my_reg[14][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat31),
	.cin(gnd),
	.combout(\my_reg[14][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[14][2]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[14][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N25
dffeas \my_reg[14][2] (
	.clk(CLK),
	.d(\my_reg[14][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[14][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[14][2] .is_wysiwyg = "true";
defparam \my_reg[14][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N27
dffeas \my_reg[15][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[15][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[15][2] .is_wysiwyg = "true";
defparam \my_reg[15][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N18
cycloneive_lcell_comb \my_reg[13][2]~feeder (
// Equation(s):
// \my_reg[13][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat31),
	.cin(gnd),
	.combout(\my_reg[13][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[13][2]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[13][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N19
dffeas \my_reg[13][2] (
	.clk(CLK),
	.d(\my_reg[13][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[13][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[13][2] .is_wysiwyg = "true";
defparam \my_reg[13][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N12
cycloneive_lcell_comb \Mux29~17 (
// Equation(s):
// \Mux29~17_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\my_reg[13][2]~q ))) # (!dcifimemload_21 & (\my_reg[12][2]~q ))))

	.dataa(\my_reg[12][2]~q ),
	.datab(\my_reg[13][2]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux29~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~17 .lut_mask = 16'hFC0A;
defparam \Mux29~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N10
cycloneive_lcell_comb \Mux29~18 (
// Equation(s):
// \Mux29~18_combout  = (dcifimemload_22 & ((\Mux29~17_combout  & ((\my_reg[15][2]~q ))) # (!\Mux29~17_combout  & (\my_reg[14][2]~q )))) # (!dcifimemload_22 & (((\Mux29~17_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[14][2]~q ),
	.datac(\my_reg[15][2]~q ),
	.datad(\Mux29~17_combout ),
	.cin(gnd),
	.combout(\Mux29~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~18 .lut_mask = 16'hF588;
defparam \Mux29~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N10
cycloneive_lcell_comb \my_reg[6][2]~feeder (
// Equation(s):
// \my_reg[6][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat31),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[6][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[6][2]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[6][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N11
dffeas \my_reg[6][2] (
	.clk(CLK),
	.d(\my_reg[6][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[6][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[6][2] .is_wysiwyg = "true";
defparam \my_reg[6][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N12
cycloneive_lcell_comb \my_reg[7][2]~feeder (
// Equation(s):
// \my_reg[7][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat31),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[7][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[7][2]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[7][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N13
dffeas \my_reg[7][2] (
	.clk(CLK),
	.d(\my_reg[7][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[7][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[7][2] .is_wysiwyg = "true";
defparam \my_reg[7][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N30
cycloneive_lcell_comb \my_reg[4][2]~feeder (
// Equation(s):
// \my_reg[4][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat31),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[4][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[4][2]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[4][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N31
dffeas \my_reg[4][2] (
	.clk(CLK),
	.d(\my_reg[4][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[4][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[4][2] .is_wysiwyg = "true";
defparam \my_reg[4][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N1
dffeas \my_reg[5][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[5][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[5][2] .is_wysiwyg = "true";
defparam \my_reg[5][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N0
cycloneive_lcell_comb \Mux29~10 (
// Equation(s):
// \Mux29~10_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\my_reg[5][2]~q ))) # (!dcifimemload_21 & (\my_reg[4][2]~q ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[4][2]~q ),
	.datac(\my_reg[5][2]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux29~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~10 .lut_mask = 16'hFA44;
defparam \Mux29~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N4
cycloneive_lcell_comb \Mux29~11 (
// Equation(s):
// \Mux29~11_combout  = (\Mux29~10_combout  & (((\my_reg[7][2]~q ) # (!dcifimemload_22)))) # (!\Mux29~10_combout  & (\my_reg[6][2]~q  & ((dcifimemload_22))))

	.dataa(\my_reg[6][2]~q ),
	.datab(\my_reg[7][2]~q ),
	.datac(\Mux29~10_combout ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux29~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~11 .lut_mask = 16'hCAF0;
defparam \Mux29~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N20
cycloneive_lcell_comb \my_reg[9][2]~feeder (
// Equation(s):
// \my_reg[9][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat31),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[9][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[9][2]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[9][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y31_N21
dffeas \my_reg[9][2] (
	.clk(CLK),
	.d(\my_reg[9][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[9][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[9][2] .is_wysiwyg = "true";
defparam \my_reg[9][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N24
cycloneive_lcell_comb \my_reg[8][2]~feeder (
// Equation(s):
// \my_reg[8][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat31),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[8][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[8][2]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[8][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N25
dffeas \my_reg[8][2] (
	.clk(CLK),
	.d(\my_reg[8][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][2] .is_wysiwyg = "true";
defparam \my_reg[8][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N2
cycloneive_lcell_comb \Mux29~12 (
// Equation(s):
// \Mux29~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][2]~q )) # (!dcifimemload_22 & ((\my_reg[8][2]~q )))))

	.dataa(\my_reg[10][2]~q ),
	.datab(\my_reg[8][2]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux29~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~12 .lut_mask = 16'hFA0C;
defparam \Mux29~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N12
cycloneive_lcell_comb \Mux29~13 (
// Equation(s):
// \Mux29~13_combout  = (dcifimemload_21 & ((\Mux29~12_combout  & (\my_reg[11][2]~q )) # (!\Mux29~12_combout  & ((\my_reg[9][2]~q ))))) # (!dcifimemload_21 & (((\Mux29~12_combout ))))

	.dataa(\my_reg[11][2]~q ),
	.datab(\my_reg[9][2]~q ),
	.datac(dcifimemload_21),
	.datad(\Mux29~12_combout ),
	.cin(gnd),
	.combout(\Mux29~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~13 .lut_mask = 16'hAFC0;
defparam \Mux29~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N16
cycloneive_lcell_comb \my_reg[3][2]~feeder (
// Equation(s):
// \my_reg[3][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat31),
	.cin(gnd),
	.combout(\my_reg[3][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[3][2]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[3][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N17
dffeas \my_reg[3][2] (
	.clk(CLK),
	.d(\my_reg[3][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[3][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[3][2] .is_wysiwyg = "true";
defparam \my_reg[3][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N2
cycloneive_lcell_comb \Mux29~14 (
// Equation(s):
// \Mux29~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][2]~q ))) # (!dcifimemload_22 & (\my_reg[1][2]~q ))))

	.dataa(\my_reg[1][2]~q ),
	.datab(\my_reg[3][2]~q ),
	.datac(dcifimemload_21),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux29~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~14 .lut_mask = 16'hC0A0;
defparam \Mux29~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N30
cycloneive_lcell_comb \my_reg[2][2]~feeder (
// Equation(s):
// \my_reg[2][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat31),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[2][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[2][2]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[2][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N31
dffeas \my_reg[2][2] (
	.clk(CLK),
	.d(\my_reg[2][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[2][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[2][2] .is_wysiwyg = "true";
defparam \my_reg[2][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N16
cycloneive_lcell_comb \Mux29~15 (
// Equation(s):
// \Mux29~15_combout  = (\Mux29~14_combout ) # ((!dcifimemload_21 & (dcifimemload_22 & \my_reg[2][2]~q )))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux29~14_combout ),
	.datad(\my_reg[2][2]~q ),
	.cin(gnd),
	.combout(\Mux29~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~15 .lut_mask = 16'hF4F0;
defparam \Mux29~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N18
cycloneive_lcell_comb \Mux29~16 (
// Equation(s):
// \Mux29~16_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\Mux29~13_combout )) # (!dcifimemload_24 & ((\Mux29~15_combout )))))

	.dataa(\Mux29~13_combout ),
	.datab(dcifimemload_23),
	.datac(dcifimemload_24),
	.datad(\Mux29~15_combout ),
	.cin(gnd),
	.combout(\Mux29~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~16 .lut_mask = 16'hE3E0;
defparam \Mux29~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N0
cycloneive_lcell_comb \my_reg[11][2]~feeder (
// Equation(s):
// \my_reg[11][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat31),
	.cin(gnd),
	.combout(\my_reg[11][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[11][2]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[11][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N1
dffeas \my_reg[11][2] (
	.clk(CLK),
	.d(\my_reg[11][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[11][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[11][2] .is_wysiwyg = "true";
defparam \my_reg[11][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N14
cycloneive_lcell_comb \Mux61~0 (
// Equation(s):
// \Mux61~0_combout  = (dcifimemload_17 & ((\my_reg[10][2]~q ) # ((dcifimemload_16)))) # (!dcifimemload_17 & (((\my_reg[8][2]~q  & !dcifimemload_16))))

	.dataa(\my_reg[10][2]~q ),
	.datab(\my_reg[8][2]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux61~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~0 .lut_mask = 16'hF0AC;
defparam \Mux61~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N8
cycloneive_lcell_comb \Mux61~1 (
// Equation(s):
// \Mux61~1_combout  = (dcifimemload_16 & ((\Mux61~0_combout  & (\my_reg[11][2]~q )) # (!\Mux61~0_combout  & ((\my_reg[9][2]~q ))))) # (!dcifimemload_16 & (((\Mux61~0_combout ))))

	.dataa(\my_reg[11][2]~q ),
	.datab(\my_reg[9][2]~q ),
	.datac(dcifimemload_16),
	.datad(\Mux61~0_combout ),
	.cin(gnd),
	.combout(\Mux61~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~1 .lut_mask = 16'hAFC0;
defparam \Mux61~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N12
cycloneive_lcell_comb \my_reg[12][2]~feeder (
// Equation(s):
// \my_reg[12][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat31),
	.cin(gnd),
	.combout(\my_reg[12][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[12][2]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[12][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N13
dffeas \my_reg[12][2] (
	.clk(CLK),
	.d(\my_reg[12][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][2] .is_wysiwyg = "true";
defparam \my_reg[12][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N24
cycloneive_lcell_comb \Mux61~7 (
// Equation(s):
// \Mux61~7_combout  = (dcifimemload_16 & ((\my_reg[13][2]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((!dcifimemload_17 & \my_reg[12][2]~q ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[13][2]~q ),
	.datac(dcifimemload_17),
	.datad(\my_reg[12][2]~q ),
	.cin(gnd),
	.combout(\Mux61~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~7 .lut_mask = 16'hADA8;
defparam \Mux61~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N26
cycloneive_lcell_comb \Mux61~8 (
// Equation(s):
// \Mux61~8_combout  = (dcifimemload_17 & ((\Mux61~7_combout  & ((\my_reg[15][2]~q ))) # (!\Mux61~7_combout  & (\my_reg[14][2]~q )))) # (!dcifimemload_17 & (((\Mux61~7_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[14][2]~q ),
	.datac(\my_reg[15][2]~q ),
	.datad(\Mux61~7_combout ),
	.cin(gnd),
	.combout(\Mux61~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~8 .lut_mask = 16'hF588;
defparam \Mux61~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N1
dffeas \my_reg[1][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[1][2] .is_wysiwyg = "true";
defparam \my_reg[1][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N0
cycloneive_lcell_comb \Mux61~4 (
// Equation(s):
// \Mux61~4_combout  = (dcifimemload_16 & ((dcifimemload_17 & (\my_reg[3][2]~q )) # (!dcifimemload_17 & ((\my_reg[1][2]~q )))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[3][2]~q ),
	.datac(\my_reg[1][2]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux61~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~4 .lut_mask = 16'h88A0;
defparam \Mux61~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N24
cycloneive_lcell_comb \Mux61~5 (
// Equation(s):
// \Mux61~5_combout  = (\Mux61~4_combout ) # ((\my_reg[2][2]~q  & (!dcifimemload_16 & dcifimemload_17)))

	.dataa(\my_reg[2][2]~q ),
	.datab(dcifimemload_16),
	.datac(\Mux61~4_combout ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux61~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~5 .lut_mask = 16'hF2F0;
defparam \Mux61~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N4
cycloneive_lcell_comb \Mux61~2 (
// Equation(s):
// \Mux61~2_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][2]~q ))) # (!dcifimemload_16 & (\my_reg[4][2]~q ))))

	.dataa(\my_reg[4][2]~q ),
	.datab(\my_reg[5][2]~q ),
	.datac(dcifimemload_17),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux61~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~2 .lut_mask = 16'hFC0A;
defparam \Mux61~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N10
cycloneive_lcell_comb \Mux61~3 (
// Equation(s):
// \Mux61~3_combout  = (dcifimemload_17 & ((\Mux61~2_combout  & (\my_reg[7][2]~q )) # (!\Mux61~2_combout  & ((\my_reg[6][2]~q ))))) # (!dcifimemload_17 & (((\Mux61~2_combout ))))

	.dataa(\my_reg[7][2]~q ),
	.datab(\my_reg[6][2]~q ),
	.datac(dcifimemload_17),
	.datad(\Mux61~2_combout ),
	.cin(gnd),
	.combout(\Mux61~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~3 .lut_mask = 16'hAFC0;
defparam \Mux61~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N18
cycloneive_lcell_comb \Mux61~6 (
// Equation(s):
// \Mux61~6_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\Mux61~3_combout ))) # (!dcifimemload_18 & (\Mux61~5_combout ))))

	.dataa(dcifimemload_19),
	.datab(\Mux61~5_combout ),
	.datac(dcifimemload_18),
	.datad(\Mux61~3_combout ),
	.cin(gnd),
	.combout(\Mux61~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~6 .lut_mask = 16'hF4A4;
defparam \Mux61~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N18
cycloneive_lcell_comb \my_reg[17][2]~feeder (
// Equation(s):
// \my_reg[17][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat31),
	.cin(gnd),
	.combout(\my_reg[17][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[17][2]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[17][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y33_N19
dffeas \my_reg[17][2] (
	.clk(CLK),
	.d(\my_reg[17][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][2] .is_wysiwyg = "true";
defparam \my_reg[17][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N2
cycloneive_lcell_comb \Mux61~10 (
// Equation(s):
// \Mux61~10_combout  = (dcifimemload_18 & ((\my_reg[21][2]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\my_reg[17][2]~q  & !dcifimemload_19))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[21][2]~q ),
	.datac(\my_reg[17][2]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux61~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~10 .lut_mask = 16'hAAD8;
defparam \Mux61~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N28
cycloneive_lcell_comb \Mux61~11 (
// Equation(s):
// \Mux61~11_combout  = (dcifimemload_19 & ((\Mux61~10_combout  & ((\my_reg[29][2]~q ))) # (!\Mux61~10_combout  & (\my_reg[25][2]~q )))) # (!dcifimemload_19 & (((\Mux61~10_combout ))))

	.dataa(\my_reg[25][2]~q ),
	.datab(\my_reg[29][2]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux61~10_combout ),
	.cin(gnd),
	.combout(\Mux61~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~11 .lut_mask = 16'hCFA0;
defparam \Mux61~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N10
cycloneive_lcell_comb \my_reg[27][2]~feeder (
// Equation(s):
// \my_reg[27][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat31),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[27][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[27][2]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[27][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N11
dffeas \my_reg[27][2] (
	.clk(CLK),
	.d(\my_reg[27][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[27][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[27][2] .is_wysiwyg = "true";
defparam \my_reg[27][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N0
cycloneive_lcell_comb \Mux61~17 (
// Equation(s):
// \Mux61~17_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & (\my_reg[23][2]~q )) # (!dcifimemload_18 & ((\my_reg[19][2]~q )))))

	.dataa(\my_reg[23][2]~q ),
	.datab(\my_reg[19][2]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux61~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~17 .lut_mask = 16'hFA0C;
defparam \Mux61~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N30
cycloneive_lcell_comb \Mux61~18 (
// Equation(s):
// \Mux61~18_combout  = (dcifimemload_19 & ((\Mux61~17_combout  & (\my_reg[31][2]~q )) # (!\Mux61~17_combout  & ((\my_reg[27][2]~q ))))) # (!dcifimemload_19 & (((\Mux61~17_combout ))))

	.dataa(\my_reg[31][2]~q ),
	.datab(\my_reg[27][2]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux61~17_combout ),
	.cin(gnd),
	.combout(\Mux61~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~18 .lut_mask = 16'hAFC0;
defparam \Mux61~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y35_N7
dffeas \my_reg[28][2] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][2] .is_wysiwyg = "true";
defparam \my_reg[28][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N20
cycloneive_lcell_comb \Mux61~14 (
// Equation(s):
// \Mux61~14_combout  = (dcifimemload_19 & ((\my_reg[24][2]~q ) # ((dcifimemload_18)))) # (!dcifimemload_19 & (((\my_reg[16][2]~q  & !dcifimemload_18))))

	.dataa(dcifimemload_19),
	.datab(\my_reg[24][2]~q ),
	.datac(\my_reg[16][2]~q ),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux61~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~14 .lut_mask = 16'hAAD8;
defparam \Mux61~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N6
cycloneive_lcell_comb \Mux61~15 (
// Equation(s):
// \Mux61~15_combout  = (dcifimemload_18 & ((\Mux61~14_combout  & ((\my_reg[28][2]~q ))) # (!\Mux61~14_combout  & (\my_reg[20][2]~q )))) # (!dcifimemload_18 & (((\Mux61~14_combout ))))

	.dataa(\my_reg[20][2]~q ),
	.datab(dcifimemload_18),
	.datac(\my_reg[28][2]~q ),
	.datad(\Mux61~14_combout ),
	.cin(gnd),
	.combout(\Mux61~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~15 .lut_mask = 16'hF388;
defparam \Mux61~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N26
cycloneive_lcell_comb \my_reg[22][2]~feeder (
// Equation(s):
// \my_reg[22][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat31),
	.cin(gnd),
	.combout(\my_reg[22][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[22][2]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[22][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y43_N27
dffeas \my_reg[22][2] (
	.clk(CLK),
	.d(\my_reg[22][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][2] .is_wysiwyg = "true";
defparam \my_reg[22][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N8
cycloneive_lcell_comb \my_reg[26][2]~feeder (
// Equation(s):
// \my_reg[26][2]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat31),
	.cin(gnd),
	.combout(\my_reg[26][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[26][2]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[26][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y43_N9
dffeas \my_reg[26][2] (
	.clk(CLK),
	.d(\my_reg[26][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][2] .is_wysiwyg = "true";
defparam \my_reg[26][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N16
cycloneive_lcell_comb \Mux61~12 (
// Equation(s):
// \Mux61~12_combout  = (dcifimemload_18 & (((dcifimemload_19)))) # (!dcifimemload_18 & ((dcifimemload_19 & (\my_reg[26][2]~q )) # (!dcifimemload_19 & ((\my_reg[18][2]~q )))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[26][2]~q ),
	.datac(\my_reg[18][2]~q ),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux61~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~12 .lut_mask = 16'hEE50;
defparam \Mux61~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N26
cycloneive_lcell_comb \Mux61~13 (
// Equation(s):
// \Mux61~13_combout  = (dcifimemload_18 & ((\Mux61~12_combout  & ((\my_reg[30][2]~q ))) # (!\Mux61~12_combout  & (\my_reg[22][2]~q )))) # (!dcifimemload_18 & (((\Mux61~12_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[22][2]~q ),
	.datac(\my_reg[30][2]~q ),
	.datad(\Mux61~12_combout ),
	.cin(gnd),
	.combout(\Mux61~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~13 .lut_mask = 16'hF588;
defparam \Mux61~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N28
cycloneive_lcell_comb \Mux61~16 (
// Equation(s):
// \Mux61~16_combout  = (dcifimemload_17 & ((dcifimemload_16) # ((\Mux61~13_combout )))) # (!dcifimemload_17 & (!dcifimemload_16 & (\Mux61~15_combout )))

	.dataa(dcifimemload_17),
	.datab(dcifimemload_16),
	.datac(\Mux61~15_combout ),
	.datad(\Mux61~13_combout ),
	.cin(gnd),
	.combout(\Mux61~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~16 .lut_mask = 16'hBA98;
defparam \Mux61~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N28
cycloneive_lcell_comb \my_reg[17][1]~feeder (
// Equation(s):
// \my_reg[17][1]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\my_reg[17][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[17][1]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[17][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N29
dffeas \my_reg[17][1] (
	.clk(CLK),
	.d(\my_reg[17][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][1] .is_wysiwyg = "true";
defparam \my_reg[17][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N16
cycloneive_lcell_comb \Mux62~0 (
// Equation(s):
// \Mux62~0_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\my_reg[25][1]~q )))) # (!dcifimemload_19 & (!dcifimemload_18 & ((\my_reg[17][1]~q ))))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\my_reg[25][1]~q ),
	.datad(\my_reg[17][1]~q ),
	.cin(gnd),
	.combout(\Mux62~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~0 .lut_mask = 16'hB9A8;
defparam \Mux62~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N30
cycloneive_lcell_comb \Mux62~1 (
// Equation(s):
// \Mux62~1_combout  = (dcifimemload_18 & ((\Mux62~0_combout  & (\my_reg[29][1]~q )) # (!\Mux62~0_combout  & ((\my_reg[21][1]~q ))))) # (!dcifimemload_18 & (((\Mux62~0_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[29][1]~q ),
	.datac(\my_reg[21][1]~q ),
	.datad(\Mux62~0_combout ),
	.cin(gnd),
	.combout(\Mux62~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~1 .lut_mask = 16'hDDA0;
defparam \Mux62~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N24
cycloneive_lcell_comb \my_reg[19][1]~feeder (
// Equation(s):
// \my_reg[19][1]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\my_reg[19][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[19][1]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[19][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y34_N25
dffeas \my_reg[19][1] (
	.clk(CLK),
	.d(\my_reg[19][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][1] .is_wysiwyg = "true";
defparam \my_reg[19][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N30
cycloneive_lcell_comb \Mux62~7 (
// Equation(s):
// \Mux62~7_combout  = (dcifimemload_19 & ((\my_reg[27][1]~q ) # ((dcifimemload_18)))) # (!dcifimemload_19 & (((\my_reg[19][1]~q  & !dcifimemload_18))))

	.dataa(\my_reg[27][1]~q ),
	.datab(\my_reg[19][1]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux62~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~7 .lut_mask = 16'hF0AC;
defparam \Mux62~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N2
cycloneive_lcell_comb \Mux62~8 (
// Equation(s):
// \Mux62~8_combout  = (dcifimemload_18 & ((\Mux62~7_combout  & ((\my_reg[31][1]~q ))) # (!\Mux62~7_combout  & (\my_reg[23][1]~q )))) # (!dcifimemload_18 & (((\Mux62~7_combout ))))

	.dataa(dcifimemload_18),
	.datab(\my_reg[23][1]~q ),
	.datac(\my_reg[31][1]~q ),
	.datad(\Mux62~7_combout ),
	.cin(gnd),
	.combout(\Mux62~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~8 .lut_mask = 16'hF588;
defparam \Mux62~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N24
cycloneive_lcell_comb \my_reg[28][1]~feeder (
// Equation(s):
// \my_reg[28][1]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat1),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[28][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[28][1]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[28][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N25
dffeas \my_reg[28][1] (
	.clk(CLK),
	.d(\my_reg[28][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][1] .is_wysiwyg = "true";
defparam \my_reg[28][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N12
cycloneive_lcell_comb \Mux62~4 (
// Equation(s):
// \Mux62~4_combout  = (dcifimemload_19 & (((dcifimemload_18)))) # (!dcifimemload_19 & ((dcifimemload_18 & ((\my_reg[20][1]~q ))) # (!dcifimemload_18 & (\my_reg[16][1]~q ))))

	.dataa(\my_reg[16][1]~q ),
	.datab(\my_reg[20][1]~q ),
	.datac(dcifimemload_19),
	.datad(dcifimemload_18),
	.cin(gnd),
	.combout(\Mux62~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~4 .lut_mask = 16'hFC0A;
defparam \Mux62~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N18
cycloneive_lcell_comb \Mux62~5 (
// Equation(s):
// \Mux62~5_combout  = (dcifimemload_19 & ((\Mux62~4_combout  & ((\my_reg[28][1]~q ))) # (!\Mux62~4_combout  & (\my_reg[24][1]~q )))) # (!dcifimemload_19 & (((\Mux62~4_combout ))))

	.dataa(\my_reg[24][1]~q ),
	.datab(\my_reg[28][1]~q ),
	.datac(dcifimemload_19),
	.datad(\Mux62~4_combout ),
	.cin(gnd),
	.combout(\Mux62~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~5 .lut_mask = 16'hCFA0;
defparam \Mux62~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y32_N5
dffeas \my_reg[26][1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[26][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[26][1] .is_wysiwyg = "true";
defparam \my_reg[26][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N24
cycloneive_lcell_comb \Mux62~2 (
// Equation(s):
// \Mux62~2_combout  = (dcifimemload_18 & ((\my_reg[22][1]~q ) # ((dcifimemload_19)))) # (!dcifimemload_18 & (((\my_reg[18][1]~q  & !dcifimemload_19))))

	.dataa(\my_reg[22][1]~q ),
	.datab(\my_reg[18][1]~q ),
	.datac(dcifimemload_18),
	.datad(dcifimemload_19),
	.cin(gnd),
	.combout(\Mux62~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~2 .lut_mask = 16'hF0AC;
defparam \Mux62~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N2
cycloneive_lcell_comb \Mux62~3 (
// Equation(s):
// \Mux62~3_combout  = (dcifimemload_19 & ((\Mux62~2_combout  & (\my_reg[30][1]~q )) # (!\Mux62~2_combout  & ((\my_reg[26][1]~q ))))) # (!dcifimemload_19 & (((\Mux62~2_combout ))))

	.dataa(\my_reg[30][1]~q ),
	.datab(dcifimemload_19),
	.datac(\my_reg[26][1]~q ),
	.datad(\Mux62~2_combout ),
	.cin(gnd),
	.combout(\Mux62~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~3 .lut_mask = 16'hBBC0;
defparam \Mux62~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N20
cycloneive_lcell_comb \Mux62~6 (
// Equation(s):
// \Mux62~6_combout  = (dcifimemload_17 & (((dcifimemload_16) # (\Mux62~3_combout )))) # (!dcifimemload_17 & (\Mux62~5_combout  & (!dcifimemload_16)))

	.dataa(dcifimemload_17),
	.datab(\Mux62~5_combout ),
	.datac(dcifimemload_16),
	.datad(\Mux62~3_combout ),
	.cin(gnd),
	.combout(\Mux62~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~6 .lut_mask = 16'hAEA4;
defparam \Mux62~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N6
cycloneive_lcell_comb \Mux62~10 (
// Equation(s):
// \Mux62~10_combout  = (dcifimemload_17 & (((dcifimemload_16)))) # (!dcifimemload_17 & ((dcifimemload_16 & ((\my_reg[5][1]~q ))) # (!dcifimemload_16 & (\my_reg[4][1]~q ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[4][1]~q ),
	.datac(\my_reg[5][1]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux62~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~10 .lut_mask = 16'hFA44;
defparam \Mux62~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N12
cycloneive_lcell_comb \Mux62~11 (
// Equation(s):
// \Mux62~11_combout  = (dcifimemload_17 & ((\Mux62~10_combout  & (\my_reg[7][1]~q )) # (!\Mux62~10_combout  & ((\my_reg[6][1]~q ))))) # (!dcifimemload_17 & (((\Mux62~10_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[7][1]~q ),
	.datac(\my_reg[6][1]~q ),
	.datad(\Mux62~10_combout ),
	.cin(gnd),
	.combout(\Mux62~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~11 .lut_mask = 16'hDDA0;
defparam \Mux62~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N24
cycloneive_lcell_comb \my_reg[12][1]~feeder (
// Equation(s):
// \my_reg[12][1]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\my_reg[12][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[12][1]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[12][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N25
dffeas \my_reg[12][1] (
	.clk(CLK),
	.d(\my_reg[12][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[12][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[12][1] .is_wysiwyg = "true";
defparam \my_reg[12][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N16
cycloneive_lcell_comb \Mux62~19 (
// Equation(s):
// \Mux62~19_combout  = (dcifimemload_16 & ((\my_reg[13][1]~q ) # ((dcifimemload_17)))) # (!dcifimemload_16 & (((\my_reg[12][1]~q  & !dcifimemload_17))))

	.dataa(\my_reg[13][1]~q ),
	.datab(\my_reg[12][1]~q ),
	.datac(dcifimemload_16),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux62~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~19 .lut_mask = 16'hF0AC;
defparam \Mux62~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N6
cycloneive_lcell_comb \Mux62~20 (
// Equation(s):
// \Mux62~20_combout  = (dcifimemload_17 & ((\Mux62~19_combout  & ((\my_reg[15][1]~q ))) # (!\Mux62~19_combout  & (\my_reg[14][1]~q )))) # (!dcifimemload_17 & (((\Mux62~19_combout ))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[14][1]~q ),
	.datac(\my_reg[15][1]~q ),
	.datad(\Mux62~19_combout ),
	.cin(gnd),
	.combout(\Mux62~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~20 .lut_mask = 16'hF588;
defparam \Mux62~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N0
cycloneive_lcell_comb \Mux62~15 (
// Equation(s):
// \Mux62~15_combout  = (ramiframload_17 & ((\my_reg[3][1]~q ))) # (!ramiframload_17 & (\my_reg[1][1]~q ))

	.dataa(gnd),
	.datab(\my_reg[1][1]~q ),
	.datac(\my_reg[3][1]~q ),
	.datad(ramiframload_17),
	.cin(gnd),
	.combout(\Mux62~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~15 .lut_mask = 16'hF0CC;
defparam \Mux62~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N18
cycloneive_lcell_comb \Mux62~16 (
// Equation(s):
// \Mux62~16_combout  = (ccifiwait_0 & (((ramiframload_16 & \Mux62~15_combout )))) # (!ccifiwait_0 & (\Mux62~14_combout ))

	.dataa(\Mux62~14_combout ),
	.datab(ccifiwait_0),
	.datac(ramiframload_16),
	.datad(\Mux62~15_combout ),
	.cin(gnd),
	.combout(\Mux62~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~16 .lut_mask = 16'hE222;
defparam \Mux62~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N14
cycloneive_lcell_comb \Mux62~17 (
// Equation(s):
// \Mux62~17_combout  = (\Mux62~16_combout ) # ((!dcifimemload_16 & (\my_reg[2][1]~q  & dcifimemload_17)))

	.dataa(dcifimemload_16),
	.datab(\Mux62~16_combout ),
	.datac(\my_reg[2][1]~q ),
	.datad(dcifimemload_17),
	.cin(gnd),
	.combout(\Mux62~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~17 .lut_mask = 16'hDCCC;
defparam \Mux62~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N16
cycloneive_lcell_comb \Mux62~12 (
// Equation(s):
// \Mux62~12_combout  = (dcifimemload_17 & ((\my_reg[10][1]~q ) # ((dcifimemload_16)))) # (!dcifimemload_17 & (((\my_reg[8][1]~q  & !dcifimemload_16))))

	.dataa(dcifimemload_17),
	.datab(\my_reg[10][1]~q ),
	.datac(\my_reg[8][1]~q ),
	.datad(dcifimemload_16),
	.cin(gnd),
	.combout(\Mux62~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~12 .lut_mask = 16'hAAD8;
defparam \Mux62~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N10
cycloneive_lcell_comb \Mux62~13 (
// Equation(s):
// \Mux62~13_combout  = (dcifimemload_16 & ((\Mux62~12_combout  & ((\my_reg[11][1]~q ))) # (!\Mux62~12_combout  & (\my_reg[9][1]~q )))) # (!dcifimemload_16 & (((\Mux62~12_combout ))))

	.dataa(dcifimemload_16),
	.datab(\my_reg[9][1]~q ),
	.datac(\my_reg[11][1]~q ),
	.datad(\Mux62~12_combout ),
	.cin(gnd),
	.combout(\Mux62~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~13 .lut_mask = 16'hF588;
defparam \Mux62~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N28
cycloneive_lcell_comb \Mux62~18 (
// Equation(s):
// \Mux62~18_combout  = (dcifimemload_19 & ((dcifimemload_18) # ((\Mux62~13_combout )))) # (!dcifimemload_19 & (!dcifimemload_18 & (\Mux62~17_combout )))

	.dataa(dcifimemload_19),
	.datab(dcifimemload_18),
	.datac(\Mux62~17_combout ),
	.datad(\Mux62~13_combout ),
	.cin(gnd),
	.combout(\Mux62~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~18 .lut_mask = 16'hBA98;
defparam \Mux62~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N4
cycloneive_lcell_comb \my_reg[22][0]~feeder (
// Equation(s):
// \my_reg[22][0]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat),
	.cin(gnd),
	.combout(\my_reg[22][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[22][0]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[22][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N5
dffeas \my_reg[22][0] (
	.clk(CLK),
	.d(\my_reg[22][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[22][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[22][0] .is_wysiwyg = "true";
defparam \my_reg[22][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N24
cycloneive_lcell_comb \Mux31~2 (
// Equation(s):
// \Mux31~2_combout  = (dcifimemload_23 & ((\my_reg[22][0]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[18][0]~q  & !dcifimemload_24))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[22][0]~q ),
	.datac(\my_reg[18][0]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~2 .lut_mask = 16'hAAD8;
defparam \Mux31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N18
cycloneive_lcell_comb \Mux31~3 (
// Equation(s):
// \Mux31~3_combout  = (dcifimemload_24 & ((\Mux31~2_combout  & ((\my_reg[30][0]~q ))) # (!\Mux31~2_combout  & (\my_reg[26][0]~q )))) # (!dcifimemload_24 & (((\Mux31~2_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[26][0]~q ),
	.datac(\my_reg[30][0]~q ),
	.datad(\Mux31~2_combout ),
	.cin(gnd),
	.combout(\Mux31~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~3 .lut_mask = 16'hF588;
defparam \Mux31~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N4
cycloneive_lcell_comb \my_reg[28][0]~feeder (
// Equation(s):
// \my_reg[28][0]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat),
	.datad(gnd),
	.cin(gnd),
	.combout(\my_reg[28][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[28][0]~feeder .lut_mask = 16'hF0F0;
defparam \my_reg[28][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N5
dffeas \my_reg[28][0] (
	.clk(CLK),
	.d(\my_reg[28][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[28][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[28][0] .is_wysiwyg = "true";
defparam \my_reg[28][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N2
cycloneive_lcell_comb \Mux31~4 (
// Equation(s):
// \Mux31~4_combout  = (dcifimemload_23 & ((\my_reg[20][0]~q ) # ((dcifimemload_24)))) # (!dcifimemload_23 & (((\my_reg[16][0]~q  & !dcifimemload_24))))

	.dataa(\my_reg[20][0]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[16][0]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux31~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~4 .lut_mask = 16'hCCB8;
defparam \Mux31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N18
cycloneive_lcell_comb \Mux31~5 (
// Equation(s):
// \Mux31~5_combout  = (dcifimemload_24 & ((\Mux31~4_combout  & (\my_reg[28][0]~q )) # (!\Mux31~4_combout  & ((\my_reg[24][0]~q ))))) # (!dcifimemload_24 & (((\Mux31~4_combout ))))

	.dataa(dcifimemload_24),
	.datab(\my_reg[28][0]~q ),
	.datac(\my_reg[24][0]~q ),
	.datad(\Mux31~4_combout ),
	.cin(gnd),
	.combout(\Mux31~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~5 .lut_mask = 16'hDDA0;
defparam \Mux31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N8
cycloneive_lcell_comb \Mux31~6 (
// Equation(s):
// \Mux31~6_combout  = (dcifimemload_21 & (dcifimemload_22)) # (!dcifimemload_21 & ((dcifimemload_22 & (\Mux31~3_combout )) # (!dcifimemload_22 & ((\Mux31~5_combout )))))

	.dataa(dcifimemload_21),
	.datab(dcifimemload_22),
	.datac(\Mux31~3_combout ),
	.datad(\Mux31~5_combout ),
	.cin(gnd),
	.combout(\Mux31~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~6 .lut_mask = 16'hD9C8;
defparam \Mux31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N5
dffeas \my_reg[17][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[17][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[17][0] .is_wysiwyg = "true";
defparam \my_reg[17][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N4
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// \Mux31~0_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[25][0]~q )) # (!dcifimemload_24 & ((\my_reg[17][0]~q )))))

	.dataa(\my_reg[25][0]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[17][0]~q ),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'hEE30;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N4
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// \Mux31~1_combout  = (dcifimemload_23 & ((\Mux31~0_combout  & ((\my_reg[29][0]~q ))) # (!\Mux31~0_combout  & (\my_reg[21][0]~q )))) # (!dcifimemload_23 & (((\Mux31~0_combout ))))

	.dataa(dcifimemload_23),
	.datab(\my_reg[21][0]~q ),
	.datac(\my_reg[29][0]~q ),
	.datad(\Mux31~0_combout ),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'hF588;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N14
cycloneive_lcell_comb \my_reg[19][0]~feeder (
// Equation(s):
// \my_reg[19][0]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat),
	.cin(gnd),
	.combout(\my_reg[19][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \my_reg[19][0]~feeder .lut_mask = 16'hFF00;
defparam \my_reg[19][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y34_N15
dffeas \my_reg[19][0] (
	.clk(CLK),
	.d(\my_reg[19][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[19][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[19][0] .is_wysiwyg = "true";
defparam \my_reg[19][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N2
cycloneive_lcell_comb \Mux31~7 (
// Equation(s):
// \Mux31~7_combout  = (dcifimemload_23 & (((dcifimemload_24)))) # (!dcifimemload_23 & ((dcifimemload_24 & (\my_reg[27][0]~q )) # (!dcifimemload_24 & ((\my_reg[19][0]~q )))))

	.dataa(\my_reg[27][0]~q ),
	.datab(\my_reg[19][0]~q ),
	.datac(dcifimemload_23),
	.datad(dcifimemload_24),
	.cin(gnd),
	.combout(\Mux31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~7 .lut_mask = 16'hFA0C;
defparam \Mux31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N20
cycloneive_lcell_comb \Mux31~8 (
// Equation(s):
// \Mux31~8_combout  = (dcifimemload_23 & ((\Mux31~7_combout  & ((\my_reg[31][0]~q ))) # (!\Mux31~7_combout  & (\my_reg[23][0]~q )))) # (!dcifimemload_23 & (((\Mux31~7_combout ))))

	.dataa(\my_reg[23][0]~q ),
	.datab(dcifimemload_23),
	.datac(\my_reg[31][0]~q ),
	.datad(\Mux31~7_combout ),
	.cin(gnd),
	.combout(\Mux31~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~8 .lut_mask = 16'hF388;
defparam \Mux31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N14
cycloneive_lcell_comb \Mux31~17 (
// Equation(s):
// \Mux31~17_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\my_reg[13][0]~q ))) # (!dcifimemload_21 & (\my_reg[12][0]~q ))))

	.dataa(\my_reg[12][0]~q ),
	.datab(dcifimemload_22),
	.datac(\my_reg[13][0]~q ),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux31~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~17 .lut_mask = 16'hFC22;
defparam \Mux31~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N0
cycloneive_lcell_comb \Mux31~18 (
// Equation(s):
// \Mux31~18_combout  = (dcifimemload_22 & ((\Mux31~17_combout  & ((\my_reg[15][0]~q ))) # (!\Mux31~17_combout  & (\my_reg[14][0]~q )))) # (!dcifimemload_22 & (((\Mux31~17_combout ))))

	.dataa(\my_reg[14][0]~q ),
	.datab(\my_reg[15][0]~q ),
	.datac(dcifimemload_22),
	.datad(\Mux31~17_combout ),
	.cin(gnd),
	.combout(\Mux31~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~18 .lut_mask = 16'hCFA0;
defparam \Mux31~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N17
dffeas \my_reg[8][0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\my_reg[8][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \my_reg[8][0] .is_wysiwyg = "true";
defparam \my_reg[8][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N16
cycloneive_lcell_comb \Mux31~12 (
// Equation(s):
// \Mux31~12_combout  = (dcifimemload_21 & (((dcifimemload_22)))) # (!dcifimemload_21 & ((dcifimemload_22 & (\my_reg[10][0]~q )) # (!dcifimemload_22 & ((\my_reg[8][0]~q )))))

	.dataa(\my_reg[10][0]~q ),
	.datab(dcifimemload_21),
	.datac(\my_reg[8][0]~q ),
	.datad(dcifimemload_22),
	.cin(gnd),
	.combout(\Mux31~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~12 .lut_mask = 16'hEE30;
defparam \Mux31~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N14
cycloneive_lcell_comb \Mux31~13 (
// Equation(s):
// \Mux31~13_combout  = (dcifimemload_21 & ((\Mux31~12_combout  & ((\my_reg[11][0]~q ))) # (!\Mux31~12_combout  & (\my_reg[9][0]~q )))) # (!dcifimemload_21 & (((\Mux31~12_combout ))))

	.dataa(dcifimemload_21),
	.datab(\my_reg[9][0]~q ),
	.datac(\my_reg[11][0]~q ),
	.datad(\Mux31~12_combout ),
	.cin(gnd),
	.combout(\Mux31~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~13 .lut_mask = 16'hF588;
defparam \Mux31~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N24
cycloneive_lcell_comb \Mux31~14 (
// Equation(s):
// \Mux31~14_combout  = (dcifimemload_21 & ((dcifimemload_22 & ((\my_reg[3][0]~q ))) # (!dcifimemload_22 & (\my_reg[1][0]~q ))))

	.dataa(\my_reg[1][0]~q ),
	.datab(\my_reg[3][0]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux31~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~14 .lut_mask = 16'hCA00;
defparam \Mux31~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N30
cycloneive_lcell_comb \Mux31~15 (
// Equation(s):
// \Mux31~15_combout  = (\Mux31~14_combout ) # ((dcifimemload_22 & (!dcifimemload_21 & \my_reg[2][0]~q )))

	.dataa(dcifimemload_22),
	.datab(dcifimemload_21),
	.datac(\my_reg[2][0]~q ),
	.datad(\Mux31~14_combout ),
	.cin(gnd),
	.combout(\Mux31~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~15 .lut_mask = 16'hFF20;
defparam \Mux31~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N22
cycloneive_lcell_comb \Mux31~16 (
// Equation(s):
// \Mux31~16_combout  = (dcifimemload_23 & (dcifimemload_24)) # (!dcifimemload_23 & ((dcifimemload_24 & (\Mux31~13_combout )) # (!dcifimemload_24 & ((\Mux31~15_combout )))))

	.dataa(dcifimemload_23),
	.datab(dcifimemload_24),
	.datac(\Mux31~13_combout ),
	.datad(\Mux31~15_combout ),
	.cin(gnd),
	.combout(\Mux31~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~16 .lut_mask = 16'hD9C8;
defparam \Mux31~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N24
cycloneive_lcell_comb \Mux31~10 (
// Equation(s):
// \Mux31~10_combout  = (dcifimemload_22 & (((dcifimemload_21)))) # (!dcifimemload_22 & ((dcifimemload_21 & ((\my_reg[5][0]~q ))) # (!dcifimemload_21 & (\my_reg[4][0]~q ))))

	.dataa(\my_reg[4][0]~q ),
	.datab(\my_reg[5][0]~q ),
	.datac(dcifimemload_22),
	.datad(dcifimemload_21),
	.cin(gnd),
	.combout(\Mux31~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~10 .lut_mask = 16'hFC0A;
defparam \Mux31~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N16
cycloneive_lcell_comb \Mux31~11 (
// Equation(s):
// \Mux31~11_combout  = (dcifimemload_22 & ((\Mux31~10_combout  & (\my_reg[7][0]~q )) # (!\Mux31~10_combout  & ((\my_reg[6][0]~q ))))) # (!dcifimemload_22 & (((\Mux31~10_combout ))))

	.dataa(dcifimemload_22),
	.datab(\my_reg[7][0]~q ),
	.datac(\my_reg[6][0]~q ),
	.datad(\Mux31~10_combout ),
	.cin(gnd),
	.combout(\Mux31~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~11 .lut_mask = 16'hDDA0;
defparam \Mux31~11 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module request_unit (
	reg_WEN1,
	reg_REN1,
	always1,
	dcifimemload_31,
	dcifimemload_29,
	Equal3,
	dcifdhit,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
output 	reg_WEN1;
output 	reg_REN1;
input 	always1;
input 	dcifimemload_31;
input 	dcifimemload_29;
input 	Equal3;
input 	dcifdhit;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \n_WEN~0_combout ;
wire \n_REN~0_combout ;


// Location: FF_X60_Y34_N9
dffeas reg_WEN(
	.clk(CLK),
	.d(\n_WEN~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(reg_WEN1),
	.prn(vcc));
// synopsys translate_off
defparam reg_WEN.is_wysiwyg = "true";
defparam reg_WEN.power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N31
dffeas reg_REN(
	.clk(CLK),
	.d(\n_REN~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(reg_REN1),
	.prn(vcc));
// synopsys translate_off
defparam reg_REN.is_wysiwyg = "true";
defparam reg_REN.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N8
cycloneive_lcell_comb \n_WEN~0 (
// Equation(s):
// \n_WEN~0_combout  = (Equal3 & (dcifimemload_31 & (!dcifdhit & dcifimemload_29)))

	.dataa(Equal3),
	.datab(dcifimemload_31),
	.datac(dcifdhit),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(\n_WEN~0_combout ),
	.cout());
// synopsys translate_off
defparam \n_WEN~0 .lut_mask = 16'h0800;
defparam \n_WEN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N30
cycloneive_lcell_comb \n_REN~0 (
// Equation(s):
// \n_REN~0_combout  = (Equal3 & (dcifimemload_31 & (!dcifdhit & !dcifimemload_29)))

	.dataa(Equal3),
	.datab(dcifimemload_31),
	.datac(dcifdhit),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(\n_REN~0_combout ),
	.cout());
// synopsys translate_off
defparam \n_REN~0 .lut_mask = 16'h0008;
defparam \n_REN~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module memory_control (
	reg_WEN,
	reg_REN,
	always1,
	ccifiwait_0,
	devpor,
	devclrn,
	devoe);
input 	reg_WEN;
input 	reg_REN;
input 	always1;
output 	ccifiwait_0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X58_Y34_N18
cycloneive_lcell_comb \ccif.iwait[0]~0 (
// Equation(s):
// ccifiwait_0 = (!reg_REN1 & (!reg_WEN1 & always1))

	.dataa(gnd),
	.datab(reg_REN),
	.datac(reg_WEN),
	.datad(always1),
	.cin(gnd),
	.combout(ccifiwait_0),
	.cout());
// synopsys translate_off
defparam \ccif.iwait[0]~0 .lut_mask = 16'h0300;
defparam \ccif.iwait[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule
