`ifndef CONTROL_UNIT_IF_VH
`define CONTROL_UNIT_IF_VH

// all types
`include "cpu_types_pkg.vh"

interface control_unit_if;
  // import types
  import cpu_types_pkg::*;

  logic      RegWEN, ALUSrc, ExtOp, zero, overflow, negative, dmemreq, imemREN, dmemwreq, halt, dhit; //imemreq to imemREN chnaged
  logic [1:0] PCSrc;
  logic [1:0] RegDest, MemtoReg;
  opcode_t  opcode;
  funct_t   funct;
  aluop_t   ALUOP;

  // control unit ports
  modport cu (
    output   dmemreq, imemREN, dmemwreq, PCSrc, RegWEN, RegDest, ExtOp, ALUSrc, ALUOP, MemtoReg, halt,
    input    zero, overflow, negative, opcode, funct, dhit
  );
  // control unit tb
  modport tb (
    input   dmemreq, imemREN, dmemwreq, PCSrc, RegWEN, RegDest, ExtOp, ALUSrc, ALUOP, MemtoReg, halt,
    output  zero, overflow, negative, opcode, funct, dhit
  );
endinterface

`endif //CONTROL_UNIT_IF_VH
