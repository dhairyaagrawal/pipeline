module control_unit (
  control_unit_if.cu cuif
);

endmodule
